LIBRARY work;
USE work.n_bit_int.ALL;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fir_filter_test is
	generic( 
		Win 			: INTEGER 	; -- Input bit width
		Wmult			: INTEGER 	;-- Multiplier bit width 2*W1
		Wadd 			: INTEGER 	;-- Adder width = Wmult+log2(L)-1
		Wout 			: INTEGER 	;-- Output bit width
		BUTTON_HIGH 	: STD_LOGIC ;
		PATTERN_SIZE	: INTEGER 	;
		RANGE_LOW 		: INTEGER 	; --pattern range: power of 2
		RANGE_HIGH 		: INTEGER 	; --must change pattern too
		LFilter  		: INTEGER 	); -- Filter length
	port (
		clk              	  : in  std_logic;
		reset                 : in  std_logic;
		o_data_buffer         : out std_logic_vector( Wout-1 downto 0);
		o_fir_coeff           : out std_logic_vector( Win-1 downto 0);
		o_input               : out std_logic_vector( Win-1 downto 0);
		read_out              : out integer );
end fir_filter_test;

architecture rtl of fir_filter_test is

	constant noisy_size : integer := 1060;
	type T_NOISY_INPUT is array(0 to noisy_size-1) of integer range RANGE_LOW to RANGE_HIGH;
	type T_COEFF_INPUT is array(0 to LFilter-1) of integer range RANGE_LOW to RANGE_HIGH;

	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--0,1,2,5,9,16,25,36,48,62,77,92,105,115,123,127,127,123,115,
	--105,92,77,62,48,36,25,16,9,5,2,1,0);

	-- L=256 RANGE -256 TO 255
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,-1,-1,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,
	--	-2,-2,-1,0,1,2,3,4,5,6,7,8,10,11,12,13,14,15,15,16,17,17,17,17,17,16,16,15,14,12,
	--	11,9,7,5,3,0,-3,-6,-9,-12,-15,-18,-21,-24,-27,-30,-33,-35,-38,-40,-42,-43,-45,-45,
	--	-46,-45,-45,-44,-42,-39,-37,-33,-29,-24,-19,-13,-7,0,8,16,24,33,42,52,62,73,83,94,
	--	105,116,127,137,148,159,169,179,188,197,206,214,221,228,234,240,244,248,251,253,255,
	--	255,253,251,248,244,240,234,228,221,214,206,197,188,179,169,159,148,137,127,116,105,
	--	94,83,73,62,52,42,33,24,16,8,0,-7,-13,-19,-24,-29,-33,-37,-39,-42,-44,-45,-45,-46,-45,
	--	-45,-43,-42,-40,-38,-35,-33,-30,-27,-24,-21,-18,-15,-12,-9,-6,-3,0,3,5,7,9,11,12,14,
	--	15,16,16,17,17,17,17,17,16,15,15,14,13,12,11,10,8,7,6,5,4,3,2,1,0,-1,-2,-2,-3,-3,-4,
	--	-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,-1,-1,0,0,0,0,0,0);

	-- L=256 RANGE -512 TO 511
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,-1,-1,-2,-2,-3,-4,-4,-5,-5,-6,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-7,-6,-5,-4,-3,
	--	-2,0,2,4,6,8,10,12,15,17,19,22,24,26,28,29,31,32,33,34,34,34,34,33,31,30,27,25,22,18,14,
	--	10,5,0,-5,-11,-17,-23,-29,-36,-42,-48,-54,-60,-66,-71,-76,-80,-84,-87,-89,-91,-91,-91,
	--	-90,-87,-84,-79,-74,-67,-58,-49,-39,-27,-14,0,15,31,48,66,85,105,125,146,167,189,210,232,
	--	254,276,298,319,339,359,378,396,414,430,445,459,471,482,491,498,504,509,511,511,509,504,
	--	498,491,482,471,459,445,430,414,396,378,359,339,319,298,276,254,232,210,189,167,146,125,
	--	105,85,66,48,31,15,0,-14,-27,-39,-49,-58,-67,-74,-79,-84,-87,-90,-91,-91,-91,-89,-87,-84,
	--	-80,-76,-71,-66,-60,-54,-48,-42,-36,-29,-23,-17,-11,-5,0,5,10,14,18,22,25,27,30,31,33,34,
	--	34,34,34,33,32,31,29,28,26,24,22,19,17,15,12,10,8,6,4,2,0,-2,-3,-4,-5,-6,-7,-8,-8,-8,-8,
	--	-8,-8,-8,-8,-7,-7,-6,-5,-5,-4,-4,-3,-2,-2,-1,-1,-1,0,0,0,0,0);

	-- L=256 RANGE -512 TO 511
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,1,0,-1,0,1,1,0,-1,-1,1,1,0,-1,-1,1,1,0,-1,-1,1,
	--	2,0,-2,-1,1,2,0,-2,-1,1,3,0,-3,-2,2,3,0,-3,-2,2,4,0,-4,-3,3,4,0,-5,-3,3,5,0,-6,-4,4,6,0,-7,-4,4,7,0,
	--	-8,-5,5,9,0,-10,-6,6,11,0,-12,-8,8,14,0,-15,-10,10,17,0,-19,-13,14,23,0,-27,-18,20,35,0,-43,-30,34,
	--	64,0,-97,-80,119,387,511,511,387,119,-80,-97,0,64,34,-30,-43,0,35,20,-18,-27,0,23,14,-13,-19,0,17,10,
	--	-10,-15,0,14,8,-8,-12,0,11,6,-6,-10,0,9,5,-5,-8,0,7,4,-4,-7,0,6,4,-4,-6,0,5,3,-3,-5,0,4,3,-3,-4,0,4,2,
	--	-2,-3,0,3,2,-2,-3,0,3,1,-1,-2,0,2,1,-1,-2,0,2,1,-1,-1,0,1,1,-1,-1,0,1,1,-1,-1,0,1,1,0,-1,0,1,0,0,-1,0,
	--	1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
	
	-- L=512 RANGE 256 TO 255
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-3,
	--	-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,
	--	-4,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,0,0,0,1,1,2,2,3,3,4,4,5,6,6,7,7,8,8,9,10,
	--	10,11,11,12,12,13,13,14,14,15,15,15,16,16,16,17,17,17,17,17,17,17,17,17,17,
	--	16,16,16,15,15,14,14,13,12,12,11,10,9,8,7,6,5,4,3,1,0,-1,-3,-4,-6,-7,-9,-10,
	--	-12,-13,-15,-16,-18,-19,-21,-23,-24,-26,-27,-29,-30,-31,-33,-34,-35,-37,-38,
	--	-39,-40,-41,-42,-43,-43,-44,-45,-45,-45,-45,-46,-46,-45,-45,-45,-44,-44,-43,
	--	-42,-41,-40,-38,-37,-35,-33,-31,-29,-27,-24,-22,-19,-16,-13,-10,-7,-4,0,4,8,
	--	11,16,20,24,28,33,38,42,47,52,57,62,67,73,78,83,89,94,99,105,110,116,121,127,
	--	132,137,143,148,153,159,164,169,174,179,184,188,193,197,202,206,210,214,218,
	--	222,225,228,231,234,237,240,242,244,246,248,250,251,252,253,254,255,255,255,
	--	255,254,253,252,251,250,248,246,244,242,240,237,234,231,228,225,222,218,214,
	--	210,206,202,197,193,188,184,179,174,169,164,159,153,148,143,137,132,127,121,
	--	116,110,105,99,94,89,83,78,73,67,62,57,52,47,42,38,33,28,24,20,16,11,8,4,0,
	--	-4,-7,-10,-13,-16,-19,-22,-24,-27,-29,-31,-33,-35,-37,-38,-40,-41,-42,-43,-44,
	--	-44,-45,-45,-45,-46,-46,-45,-45,-45,-45,-44,-43,-43,-42,-41,-40,-39,-38,-37,
	--	-35,-34,-33,-31,-30,-29,-27,-26,-24,-23,-21,-19,-18,-16,-15,-13,-12,-10,-9,-7,
	--	-6,-4,-3,-1,0,1,3,4,5,6,7,8,9,10,11,12,12,13,14,14,15,15,16,16,16,17,17,17,17,
	--	17,17,17,17,17,17,16,16,16,15,15,15,14,14,13,13,12,12,11,11,10,10,9,8,8,7,7,6,
	--	6,5,4,4,3,3,2,2,1,1,0,0,0,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,
	--	-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-1,-1,
	--	-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0);

	-- L=512 RANGE -512 TO 511 (1)
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,0,0,-1,-1,-1,-2,-2,-1,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,0,1,1,2,3,3,3,2,1,0,-1,-2,-3,-3,-3,-3,-3,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-4,-5,-5,-5,-4,-3,-1,1,2,4,5,6,6,5,3,2,-1,-3,-5,-6,-7,-7,-6,-4,-2,0,3,5,7,8,8,7,5,3,0,-3,-6,-8,-9,-9,-8,-6,-3,0,4,7,9,11,11,10,8,4,0,-4,-8,-11,-13,-13,-12,-9,-6,-1,4,9,12,15,15,14,11,7,2,-4,-10,-14,-17,-18,-17,-14,-9,-3,4,11,17,21,22,21,17,11,4,-5,-13,-20,-25,-27,-26,-22,-15,-6,5,15,24,31,34,33,28,20,8,-5,-18,-30,-40,-45,-44,-39,-28,-13,5,24,41,55,63,64,57,43,21,-5,-34,-63,-87,-104,-110,-104,-82,-46,5,68,139,216,292,363,424,471,501,511,511,501,471,424,363,292,216,139,68,5,-46,-82,-104,-110,-104,-87,-63,-34,-5,21,43,57,64,63,55,41,24,5,-13,-28,-39,-44,-45,-40,-30,-18,-5,8,20,28,33,34,31,24,15,5,-6,-15,-22,-26,-27,-25,-20,-13,-5,4,11,17,21,22,21,17,11,4,-3,-9,-14,-17,-18,-17,-14,-10,-4,2,7,11,14,15,15,12,9,4,-1,-6,-9,-12,-13,-13,-11,-8,-4,0,4,8,10,11,11,9,7,4,0,-3,-6,-8,-9,-9,-8,-6,-3,0,3,5,7,8,8,7,5,3,0,-2,-4,-6,-7,-7,-6,-5,-3,-1,2,3,5,6,6,5,4,2,1,-1,-3,-4,-5,-5,-5,-4,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-3,-3,-3,-3,-3,-2,-1,0,1,2,3,3,3,2,1,1,0,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-1,-2,-2,-1,-1,-1,0,0,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,-1,0,0,0,0,0
	--);
	
    -- L=512 RANGE -512 TO 511 SEM JANELA
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	4,3,1,-1,-3,-4,-4,-4,-3,-1,1,3,4,4,4,2,0,-2,-4,-5,-4,-3,-1,1,3,4,5,4,3,1,-1,-3,-5,-5,-4,-2,0,2,4,5,5,4,2,-1,-3,-5,-5,-5,-3,-1,2,4,5,5,4,2,0,-2,-4,-5,-5,-4,-2,1,3,5,6,5,3,1,-2,-4,-6,-6,-5,-3,0,3,5,6,6,4,2,-1,-4,-6,-6,-6,-4,-1,2,5,6,7,5,3,0,-3,-6,-7,-7,-5,-2,1,4,6,7,6,4,1,-2,-5,-7,-7,-6,-3,0,4,6,8,8,6,3,-1,-5,-7,-8,-7,-5,-1,3,6,8,9,7,4,0,-4,-7,-9,-9,-7,-3,2,6,9,10,9,6,2,-3,-7,-10,-10,-9,-5,0,5,9,11,11,8,4,-2,-7,-11,-12,-11,-7,-2,4,9,12,13,11,6,0,-6,-11,-14,-14,-10,-5,2,9,14,15,14,9,3,-5,-12,-16,-17,-14,-8,0,8,15,19,18,14,6,-3,-12,-19,-22,-20,-13,-4,7,17,23,25,21,12,0,-13,-23,-29,-29,-22,-10,5,20,31,36,33,23,6,-13,-31,-43,-47,-40,-23,0,26,49,63,64,51,24,-13,-53,-88,-108,-107,-80,-24,56,153,258,357,439,492,511,492,439,357,258,153,56,-24,-80,-107,-108,-88,-53,-13,24,51,64,63,49,26,0,-23,-40,-47,-43,-31,-13,6,23,33,36,31,20,5,-10,-22,-29,-29,-23,-13,0,12,21,25,23,17,7,-4,-13,-20,-22,-19,-12,-3,6,14,18,19,15,8,0,-8,-14,-17,-16,-12,-5,3,9,14,15,14,9,2,-5,-10,-14,-14,-11,-6,0,6,11,13,12,9,4,-2,-7,-11,-12,-11,-7,-2,4,8,11,11,9,5,0,-5,-9,-10,-10,-7,-3,2,6,9,10,9,6,2,-3,-7,-9,-9,-7,-4,0,4,7,9,8,6,3,-1,-5,-7,-8,-7,-5,-1,3,6,8,8,6,4,0,-3,-6,-7,-7,-5,-2,1,4,6,7,6,4,1,-2,-5,-7,-7,-6,-3,0,3,5,7,6,5,2,-1,-4,-6,-6,-6,-4,-1,2,4,6,6,5,3,0,-3,-5,-6,-6,-4,-2,1,3,5,6,5,3,1,-2,-4,-5,-5,-4,-2,0,2,4,5,5,4,2,-1,-3,-5,-5,-5,-3,-1,2,4,5,5,4,2,0,-2,-4,-5,-5,-3,-1,1,3,4,5,4,3,1,-1,-3,-4,-5,-4,-2,0,2,4,4,4,3,1,-1,-3,-4,-4,-4,-3,-1,1,3
	--);	
	
	-- L=512 RANGE -512 TO 511 (hamming) b=0.15
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,0,0,-1,-1,-1,-2,-2,-1,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,0,1,1,2,3,3,3,2,1,0,-1,-2,-3,-3,-3,-3,-3,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-4,-5,-5,-5,-4,-3,-1,1,2,4,5,6,6,5,3,2,-1,-3,-5,-6,-7,-7,-6,-4,-2,0,3,5,7,8,8,7,5,3,0,-3,-6,-8,-9,-9,-8,-6,-3,0,4,7,9,11,11,10,8,4,0,-4,-8,-11,-13,-13,-12,-9,-6,-1,4,9,12,15,15,14,11,7,2,-4,-10,-14,-17,-18,-17,-14,-9,-3,4,11,17,21,22,21,17,11,4,-5,-13,-20,-25,-27,-26,-22,-15,-6,5,15,24,31,34,33,28,20,8,-5,-18,-30,-40,-45,-44,-39,-28,-13,5,24,41,55,63,64,57,43,21,-5,-34,-63,-87,-104,-110,-104,-82,-46,5,68,139,216,292,363,424,471,501,511,511,501,471,424,363,292,216,139,68,5,-46,-82,-104,-110,-104,-87,-63,-34,-5,21,43,57,64,63,55,41,24,5,-13,-28,-39,-44,-45,-40,-30,-18,-5,8,20,28,33,34,31,24,15,5,-6,-15,-22,-26,-27,-25,-20,-13,-5,4,11,17,21,22,21,17,11,4,-3,-9,-14,-17,-18,-17,-14,-10,-4,2,7,11,14,15,15,12,9,4,-1,-6,-9,-12,-13,-13,-11,-8,-4,0,4,8,10,11,11,9,7,4,0,-3,-6,-8,-9,-9,-8,-6,-3,0,3,5,7,8,8,7,5,3,0,-2,-4,-6,-7,-7,-6,-5,-3,-1,2,3,5,6,6,5,4,2,1,-1,-3,-4,-5,-5,-5,-4,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-3,-3,-3,-3,-3,-2,-1,0,1,2,3,3,3,2,1,1,0,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-1,-2,-2,-1,-1,-1,0,0,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,-1,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (hamming) b=0.05
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,1,1,1,0,0,-1,-1,-2,-2,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-2,-2,-1,0,0,1,2,3,3,4,5,5,5,6,6,6,5,5,4,4,3,2,1,0,-2,-3,-4,-5,-6,-7,-8,-9,-9,-9,-9,-9,-9,-8,-7,-6,-5,-4,-2,0,1,3,5,7,8,10,11,12,12,13,13,13,12,11,10,8,6,4,2,0,-3,-5,-8,-10,-13,-15,-16,-18,-19,-19,-19,-19,-18,-17,-15,-13,-10,-7,-4,0,3,7,10,14,17,20,22,24,26,27,27,26,25,23,21,17,14,9,5,0,-6,-11,-16,-21,-25,-30,-33,-36,-38,-39,-40,-39,-37,-35,-31,-26,-21,-15,-8,0,7,15,23,30,37,44,49,54,57,59,60,59,57,53,47,40,32,22,11,0,-13,-26,-38,-51,-63,-75,-85,-94,-101,-106,-108,-108,-105,-99,-90,-79,-63,-45,-24,0,26,55,86,118,152,187,221,256,291,324,356,386,413,438,460,478,492,503,509,511,511,509,503,492,478,460,438,413,386,356,324,291,256,221,187,152,118,86,55,26,0,-24,-45,-63,-79,-90,-99,-105,-108,-108,-106,-101,-94,-85,-75,-63,-51,-38,-26,-13,0,11,22,32,40,47,53,57,59,60,59,57,54,49,44,37,30,23,15,7,0,-8,-15,-21,-26,-31,-35,-37,-39,-40,-39,-38,-36,-33,-30,-25,-21,-16,-11,-6,0,5,9,14,17,21,23,25,26,27,27,26,24,22,20,17,14,10,7,3,0,-4,-7,-10,-13,-15,-17,-18,-19,-19,-19,-19,-18,-16,-15,-13,-10,-8,-5,-3,0,2,4,6,8,10,11,12,13,13,13,12,12,11,10,8,7,5,3,1,0,-2,-4,-5,-6,-7,-8,-9,-9,-9,-9,-9,-9,-8,-7,-6,-5,-4,-3,-2,0,1,2,3,4,4,5,5,6,6,6,5,5,5,4,3,3,2,1,0,0,-1,-2,-2,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-2,-2,-1,-1,0,0,1,1,1,2,2,2,2,2,2,2,2,2,1,1,1,1,0,0,0,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0
	--);
	
	-- L=512 RANGE -512 TO 511 (hamming) b=0.01
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-5,-5,-6,-6,-7,-7,-8,-9,-9,-10,-11,-11,-12,-13,-14,-14,-15,-16,-17,-18,-19,-20,-21,-22,-23,-24,-25,-26,-27,-28,-29,-30,-31,-32,-33,-34,-35,-37,-38,-39,-40,-41,-42,-43,-44,-45,-46,-47,-48,-49,-50,-51,-52,-53,-54,-54,-55,-56,-57,-57,-58,-58,-59,-59,-59,-60,-60,-60,-60,-60,-60,-59,-59,-59,-58,-58,-57,-56,-56,-55,-54,-52,-51,-50,-48,-47,-45,-43,-41,-39,-37,-35,-33,-30,-27,-25,-22,-19,-16,-12,-9,-5,-2,2,6,10,14,18,23,27,32,37,42,47,52,57,62,68,73,79,85,91,97,103,109,115,121,128,134,141,148,154,161,168,175,182,189,196,203,210,217,224,231,238,246,253,260,267,274,282,289,296,303,310,317,324,331,338,344,351,358,364,371,377,383,390,396,402,407,413,419,424,430,435,440,445,450,454,459,463,467,471,475,478,482,485,488,491,494,496,499,501,503,504,506,507,508,509,510,511,511,511,511,510,509,508,507,506,504,503,501,499,496,494,491,488,485,482,478,475,471,467,463,459,454,450,445,440,435,430,424,419,413,407,402,396,390,383,377,371,364,358,351,344,338,331,324,317,310,303,296,289,282,274,267,260,253,246,238,231,224,217,210,203,196,189,182,175,168,161,154,148,141,134,128,121,115,109,103,97,91,85,79,73,68,62,57,52,47,42,37,32,27,23,18,14,10,6,2,-2,-5,-9,-12,-16,-19,-22,-25,-27,-30,-33,-35,-37,-39,-41,-43,-45,-47,-48,-50,-51,-52,-54,-55,-56,-56,-57,-58,-58,-59,-59,-59,-60,-60,-60,-60,-60,-60,-59,-59,-59,-58,-58,-57,-57,-56,-55,-54,-54,-53,-52,-51,-50,-49,-48,-47,-46,-45,-44,-43,-42,-41,-40,-39,-38,-37,-35,-34,-33,-32,-31,-30,-29,-28,-27,-26,-25,-24,-23,-22,-21,-20,-19,-18,-17,-16,-15,-14,-14,-13,-12,-11,-11,-10,-9,-9,-8,-7,-7,-6,-6,-5,-5,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.1
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,3,3,3,2,2,1,0,-1,-2,-3,-3,-4,-4,-3,-2,-1,0,1,3,4,4,5,5,4,3,2,0,-2,-3,-5,-6,-6,-6,-5,-4,-2,0,2,4,6,7,8,7,6,5,3,0,-3,-5,-7,-9,-10,-9,-8,-6,-3,0,3,7,9,11,12,12,10,8,4,0,-4,-8,-12,-14,-15,-15,-13,-10,-5,0,5,11,15,18,19,19,16,12,7,0,-7,-13,-19,-23,-24,-24,-21,-16,-8,0,9,17,24,29,32,31,27,20,11,0,-12,-23,-33,-40,-43,-42,-37,-28,-15,0,16,33,47,57,63,62,55,42,23,0,-26,-52,-76,-95,-107,-109,-100,-79,-45,0,56,119,187,257,325,386,438,478,503,511,511,503,478,438,386,325,257,187,119,56,0,-45,-79,-100,-109,-107,-95,-76,-52,-26,0,23,42,55,62,63,57,47,33,16,0,-15,-28,-37,-42,-43,-40,-33,-23,-12,0,11,20,27,31,32,29,24,17,9,0,-8,-16,-21,-24,-24,-23,-19,-13,-7,0,7,12,16,19,19,18,15,11,5,0,-5,-10,-13,-15,-15,-14,-12,-8,-4,0,4,8,10,12,12,11,9,7,3,0,-3,-6,-8,-9,-10,-9,-7,-5,-3,0,3,5,6,7,8,7,6,4,2,0,-2,-4,-5,-6,-6,-6,-5,-3,-2,0,2,3,4,5,5,4,4,3,1,0,-1,-2,-3,-4,-4,-3,-3,-2,-1,0,1,2,2,3,3,3,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	
	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.05
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,2,2,2,2,2,3,3,3,2,2,2,2,1,1,1,0,-1,-1,-2,-2,-3,-3,-4,-4,-5,-5,-5,-5,-5,-4,-4,-3,-3,-2,-1,0,1,2,3,4,5,6,7,7,8,8,8,8,8,7,7,6,4,3,2,0,-2,-3,-5,-7,-8,-10,-11,-12,-13,-14,-14,-13,-13,-12,-11,-9,-7,-5,-3,0,3,6,8,11,14,16,18,20,21,22,22,21,21,19,17,15,12,8,4,0,-4,-9,-13,-17,-22,-25,-28,-31,-33,-34,-35,-34,-33,-30,-27,-23,-18,-13,-7,0,7,14,21,28,35,41,46,50,54,56,56,56,54,50,45,39,31,21,11,0,-12,-24,-37,-49,-61,-72,-82,-91,-98,-103,-105,-105,-103,-97,-89,-77,-62,-44,-24,0,26,55,85,118,151,186,221,256,290,323,355,385,413,438,459,478,492,503,509,511,511,509,503,492,478,459,438,413,385,355,323,290,256,221,186,151,118,85,55,26,0,-24,-44,-62,-77,-89,-97,-103,-105,-105,-103,-98,-91,-82,-72,-61,-49,-37,-24,-12,0,11,21,31,39,45,50,54,56,56,56,54,50,46,41,35,28,21,14,7,0,-7,-13,-18,-23,-27,-30,-33,-34,-35,-34,-33,-31,-28,-25,-22,-17,-13,-9,-4,0,4,8,12,15,17,19,21,21,22,22,21,20,18,16,14,11,8,6,3,0,-3,-5,-7,-9,-11,-12,-13,-13,-14,-14,-13,-12,-11,-10,-8,-7,-5,-3,-2,0,2,3,4,6,7,7,8,8,8,8,8,7,7,6,5,4,3,2,1,0,-1,-2,-3,-3,-4,-4,-5,-5,-5,-5,-5,-4,-4,-3,-3,-2,-2,-1,-1,0,1,1,1,2,2,2,2,3,3,3,2,2,2,2,2,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.01
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-4,-4,-5,-5,-5,-6,-6,-7,-7,-8,-8,-9,-9,-10,-10,-11,-11,-12,-12,-13,-14,-14,-15,-16,-16,-17,-18,-18,-19,-20,-21,-21,-22,-23,-23,-24,-25,-25,-26,-27,-27,-28,-29,-29,-30,-30,-31,-31,-32,-32,-32,-33,-33,-33,-34,-34,-34,-34,-34,-34,-33,-33,-33,-33,-32,-32,-31,-30,-29,-29,-28,-27,-25,-24,-23,-21,-20,-18,-16,-14,-12,-10,-8,-6,-3,0,2,5,8,11,15,18,22,25,29,33,37,41,46,50,55,59,64,69,74,79,85,90,96,101,107,113,119,125,131,138,144,151,157,164,171,178,184,191,198,206,213,220,227,234,242,249,256,264,271,278,286,293,300,307,315,322,329,336,343,350,357,364,370,377,384,390,396,403,409,415,421,426,432,437,443,448,453,457,462,466,471,475,478,482,485,489,492,495,497,500,502,504,505,507,508,509,510,511,511,511,511,510,509,508,507,505,504,502,500,497,495,492,489,485,482,478,475,471,466,462,457,453,448,443,437,432,426,421,415,409,403,396,390,384,377,370,364,357,350,343,336,329,322,315,307,300,293,286,278,271,264,256,249,242,234,227,220,213,206,198,191,184,178,171,164,157,151,144,138,131,125,119,113,107,101,96,90,85,79,74,69,64,59,55,50,46,41,37,33,29,25,22,18,15,11,8,5,2,0,-3,-6,-8,-10,-12,-14,-16,-18,-20,-21,-23,-24,-25,-27,-28,-29,-29,-30,-31,-32,-32,-33,-33,-33,-33,-34,-34,-34,-34,-34,-34,-33,-33,-33,-32,-32,-32,-31,-31,-30,-30,-29,-29,-28,-27,-27,-26,-25,-25,-24,-23,-23,-22,-21,-21,-20,-19,-18,-18,-17,-16,-16,-15,-14,-14,-13,-12,-12,-11,-11,-10,-10,-9,-9,-8,-8,-7,-7,-6,-6,-5,-5,-5,-4,-4,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 ofdm hamming
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,-1,0,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-2,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-2,2,0,-3,1,2,-2,-1,3,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-4,1,3,-3,-2,4,-1,-4,3,2,-5,0,5,-3,-3,5,0,-5,3,4,-6,0,6,-3,-4,6,1,-7,3,6,-7,-2,8,-3,-7,8,3,-10,4,9,-9,-4,13,-4,-12,11,6,-17,4,17,-15,-10,24,-4,-27,23,20,-44,4,64,-56,-77,261,511,261,-77,-56,64,4,-44,20,23,-27,-4,24,-10,-15,17,4,-17,6,11,-12,-4,13,-4,-9,9,4,-10,3,8,-7,-3,8,-2,-7,6,3,-7,1,6,-4,-3,6,0,-6,4,3,-5,0,5,-3,-3,5,0,-5,2,3,-4,-1,4,-2,-3,3,1,-4,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,3,-1,-2,2,1,-3,0,2,-2,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,1,0,-2,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,0,-1,0,1,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);

	-- >>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>JANELAS
	-- L=512 RANGE -1024 TO 1023 ofdm hamming 1
	constant COEFF_ARRAY : T_COEFF_INPUT := (
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-3,1,2,-2,-1,3,-1,-3,2,1,-3,1,3,-2,-1,3,-1,-3,3,2,-4,0,4,-3,-2,4,0,-4,3,3,-4,0,5,-2,-3,5,1,-5,2,4,-5,-1,6,-2,-4,5,2,-6,2,5,-5,-2,7,-2,-6,6,3,-8,2,7,-6,-4,8,-1,-8,6,5,-9,1,9,-6,-6,10,0,-11,6,7,-11,-1,12,-7,-9,12,2,-14,7,11,-14,-3,17,-7,-14,16,5,-21,7,18,-19,-8,26,-7,-24,23,12,-34,7,34,-30,-20,49,-7,-55,46,40,-89,7,127,-113,-155,522,1023,522,-155,-113,127,7,-89,40,46,-55,-7,49,-20,-30,34,7,-34,12,23,-24,-7,26,-8,-19,18,7,-21,5,16,-14,-7,17,-3,-14,11,7,-14,2,12,-9,-7,12,-1,-11,7,6,-11,0,10,-6,-6,9,1,-9,5,6,-8,-1,8,-4,-6,7,2,-8,3,6,-6,-2,7,-2,-5,5,2,-6,2,5,-4,-2,6,-1,-5,4,2,-5,1,5,-3,-2,5,0,-4,3,3,-4,0,4,-2,-3,4,0,-4,2,3,-3,-1,3,-1,-2,3,1,-3,1,2,-3,-1,3,-1,-2,2,1,-3,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);
	-- L=512 RANGE -1024 TO 1023 ofdm blackman 2
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,2,-1,-1,1,0,-2,1,1,-2,-1,2,-1,-2,2,1,-2,0,2,-2,-1,3,0,-2,2,1,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,4,-2,-3,4,1,-4,2,3,-4,-1,5,-2,-4,4,1,-5,2,4,-5,-2,6,-2,-5,5,3,-7,1,6,-5,-3,8,-1,-7,6,4,-8,1,8,-6,-5,9,0,-10,6,7,-11,-1,12,-6,-9,12,2,-14,7,11,-14,-3,17,-7,-14,16,5,-20,7,18,-19,-8,25,-7,-24,23,12,-33,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-33,12,23,-24,-7,25,-8,-19,18,7,-20,5,16,-14,-7,17,-3,-14,11,7,-14,2,12,-9,-6,12,-1,-11,7,6,-10,0,9,-5,-6,8,1,-8,4,6,-7,-1,8,-3,-5,6,1,-7,3,5,-5,-2,6,-2,-5,4,2,-5,1,4,-4,-2,5,-1,-4,3,2,-4,1,4,-3,-2,4,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,1,2,-2,0,3,-1,-2,2,0,-2,1,2,-2,-1,2,-1,-2,1,1,-2,0,1,-1,-1,2,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);	
	-- L=512 RANGE -1024 TO 1023 ofdm kaiser 3
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	-1,-2,2,1,-2,1,2,-1,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,2,-2,-1,3,0,-2,2,1,-3,0,3,-2,-1,3,0,-3,2,2,-3,0,3,-1,-2,3,0,-3,1,2,-3,0,3,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,4,0,-3,3,2,-3,0,3,-2,-2,4,0,-4,2,2,-4,0,4,-2,-3,4,1,-4,2,3,-4,-1,4,-2,-3,4,1,-4,2,4,-4,-1,5,-1,-4,4,2,-5,1,4,-4,-2,5,-1,-5,4,3,-5,1,5,-3,-3,6,0,-5,3,4,-6,0,6,-3,-4,6,1,-6,3,5,-6,-1,7,-3,-5,6,2,-7,3,6,-6,-2,8,-2,-7,7,3,-9,2,8,-7,-4,9,-1,-9,7,5,-10,1,10,-7,-6,11,0,-11,7,8,-12,-1,13,-7,-9,13,2,-15,7,12,-14,-3,18,-7,-14,17,5,-21,7,18,-19,-8,26,-7,-24,23,13,-34,7,34,-30,-20,49,-7,-55,46,40,-89,7,128,-113,-155,522,1023,522,-155,-113,128,7,-89,40,46,-55,-7,49,-20,-30,34,7,-34,13,23,-24,-7,26,-8,-19,18,7,-21,5,17,-14,-7,18,-3,-14,12,7,-15,2,13,-9,-7,13,-1,-12,8,7,-11,0,11,-6,-7,10,1,-10,5,7,-9,-1,9,-4,-7,8,2,-9,3,7,-7,-2,8,-2,-6,6,3,-7,2,6,-5,-3,7,-1,-6,5,3,-6,1,6,-4,-3,6,0,-6,4,3,-5,0,6,-3,-3,5,1,-5,3,4,-5,-1,5,-2,-4,4,1,-5,2,4,-4,-1,5,-1,-4,4,2,-4,1,4,-3,-2,4,-1,-4,3,2,-4,1,4,-3,-2,4,0,-4,2,2,-4,0,4,-2,-2,3,0,-3,2,3,-3,0,4,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,3,0,-3,2,1,-3,0,3,-2,-1,3,0,-3,2,2,-3,0,3,-1,-2,3,0,-3,1,2,-2,0,3,-1,-2,2,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-1,2,1,-2,1,2,-2,-1,2
	--);
	-- L=512 RANGE -1024 TO 1023 ofdm Chebyshev 4
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,2,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,2,1,-2,0,2,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-4,2,3,-4,-1,4,-2,-3,4,1,-5,2,4,-4,-2,5,-2,-5,5,2,-6,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-6,-5,9,0,-10,6,7,-10,-1,11,-6,-8,12,2,-13,6,10,-13,-3,16,-7,-13,15,5,-20,7,17,-18,-8,25,-7,-24,23,12,-33,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-33,12,23,-24,-7,25,-8,-18,17,7,-20,5,15,-13,-7,16,-3,-13,10,6,-13,2,12,-8,-6,11,-1,-10,7,6,-10,0,9,-5,-6,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-6,2,5,-5,-2,5,-2,-4,4,2,-5,1,4,-3,-2,4,-1,-4,3,2,-4,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,2,0,-2,1,2,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,2,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- L=512 RANGE -1024 TO 1023 ofdm Barltlett-Hann 5
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,4,0,-4,2,3,-4,0,4,-2,-3,4,1,-5,2,4,-5,-1,5,-2,-4,5,1,-6,2,5,-5,-2,7,-2,-6,5,3,-7,2,7,-6,-3,8,-1,-8,6,4,-9,1,9,-6,-6,10,0,-10,6,7,-11,-1,12,-6,-9,12,2,-14,7,11,-14,-3,17,-7,-14,16,5,-20,7,18,-18,-8,25,-7,-24,23,12,-33,7,34,-30,-20,48,-7,-54,45,39,-88,7,127,-113,-154,522,1023,522,-154,-113,127,7,-88,39,45,-54,-7,48,-20,-30,34,7,-33,12,23,-24,-7,25,-8,-18,18,7,-20,5,16,-14,-7,17,-3,-14,11,7,-14,2,12,-9,-6,12,-1,-11,7,6,-10,0,10,-6,-6,9,1,-9,4,6,-8,-1,8,-3,-6,7,2,-7,3,5,-6,-2,7,-2,-5,5,2,-6,1,5,-4,-2,5,-1,-5,4,2,-5,1,4,-3,-2,4,0,-4,3,2,-4,0,4,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Barltlett 6
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-4,2,2,-4,0,4,-2,-3,4,1,-4,2,3,-4,-1,5,-2,-4,4,1,-5,2,4,-5,-2,6,-2,-5,5,2,-7,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-5,-5,9,0,-9,6,6,-10,-1,11,-6,-8,11,2,-13,6,10,-13,-3,15,-6,-13,15,5,-19,7,17,-17,-7,24,-7,-22,22,12,-32,7,32,-29,-20,47,-7,-53,44,39,-87,7,126,-112,-153,520,1023,520,-153,-112,126,7,-87,39,44,-53,-7,47,-20,-29,32,7,-32,12,22,-22,-7,24,-7,-17,17,7,-19,5,15,-13,-6,15,-3,-13,10,6,-13,2,11,-8,-6,11,-1,-10,6,6,-9,0,9,-5,-5,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-7,2,5,-5,-2,6,-2,-5,4,2,-5,1,4,-4,-2,5,-1,-4,3,2,-4,1,4,-3,-2,4,0,-4,2,2,-4,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Blackman-Harris 7
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-2,-1,2,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,2,3,-3,-1,4,-2,-3,4,1,-5,2,4,-4,-2,5,-1,-5,4,2,-6,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-5,-5,9,0,-9,6,6,-10,-1,11,-6,-8,12,2,-13,6,10,-13,-3,16,-7,-13,15,5,-20,7,17,-18,-8,25,-7,-23,23,12,-33,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-33,12,23,-23,-7,25,-8,-18,17,7,-20,5,15,-13,-7,16,-3,-13,10,6,-13,2,12,-8,-6,11,-1,-10,6,6,-9,0,9,-5,-5,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-6,2,4,-5,-1,5,-2,-4,4,2,-5,1,4,-3,-2,4,-1,-3,3,2,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,2,-1,-2,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- L=512 RANGE -1024 TO 1023 ofdm Bohman 8
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-2,1,1,-1,-1,2,-1,-2,2,1,-2,0,2,-2,-1,2,0,-2,2,1,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,4,-2,-3,4,0,-4,2,3,-4,-1,5,-2,-4,4,1,-5,2,4,-5,-2,6,-2,-5,5,2,-7,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-6,-5,9,0,-10,6,7,-10,-1,12,-6,-8,12,2,-14,7,11,-13,-3,16,-7,-14,16,5,-20,7,18,-18,-8,25,-7,-24,23,12,-33,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-33,12,23,-24,-7,25,-8,-18,18,7,-20,5,16,-14,-7,16,-3,-13,11,7,-14,2,12,-8,-6,12,-1,-10,7,6,-10,0,9,-5,-6,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-7,2,5,-5,-2,6,-2,-5,4,2,-5,1,4,-4,-2,5,-1,-4,3,2,-4,0,4,-3,-2,4,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,1,2,-2,0,2,-1,-2,2,0,-2,1,2,-2,-1,2,-1,-1,1,1,-2,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Flat Top 9
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,1,-1,0,1,-1,-1,1,0,-1,1,1,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-3,3,1,-4,1,4,-3,-2,5,-1,-5,4,3,-6,0,6,-4,-4,7,0,-8,5,5,-8,-1,9,-5,-7,10,1,-12,6,9,-12,-3,15,-6,-12,14,5,-19,6,16,-17,-7,24,-7,-23,22,12,-32,7,33,-29,-20,48,-7,-54,45,39,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,39,45,-54,-7,48,-20,-29,33,7,-32,12,22,-23,-7,24,-7,-17,16,6,-19,5,14,-12,-6,15,-3,-12,9,6,-12,1,10,-7,-5,9,-1,-8,5,5,-8,0,7,-4,-4,6,0,-6,3,4,-5,-1,5,-2,-3,4,1,-4,1,3,-3,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,1,1,-1,0,1,-1,-1,1,0,-1,1,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Gaussiana 10
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,4,0,-4,2,2,-4,0,4,-2,-3,4,1,-5,2,4,-4,-1,5,-2,-4,5,1,-6,2,5,-5,-2,6,-2,-6,5,3,-7,2,7,-6,-3,8,-1,-8,6,4,-9,1,9,-6,-6,10,0,-10,6,7,-11,-1,12,-7,-9,12,2,-14,7,11,-14,-3,17,-7,-14,16,5,-20,7,18,-19,-8,25,-7,-24,23,12,-34,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-34,12,23,-24,-7,25,-8,-19,18,7,-20,5,16,-14,-7,17,-3,-14,11,7,-14,2,12,-9,-7,12,-1,-11,7,6,-10,0,10,-6,-6,9,1,-9,4,6,-8,-1,8,-3,-6,7,2,-7,3,5,-6,-2,6,-2,-5,5,2,-6,1,5,-4,-2,5,-1,-4,4,2,-5,1,4,-3,-2,4,0,-4,2,2,-4,0,4,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Hann 11
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,0,-3,2,2,-4,0,4,-2,-2,4,0,-4,2,3,-4,0,4,-2,-3,4,1,-5,2,4,-5,-1,5,-2,-4,5,2,-6,2,5,-5,-2,7,-2,-6,5,3,-7,2,7,-6,-4,8,-1,-8,6,5,-9,1,9,-6,-6,10,0,-10,6,7,-11,-1,12,-7,-9,12,2,-14,7,11,-14,-3,17,-7,-14,16,5,-20,7,18,-19,-8,26,-7,-24,23,12,-34,7,34,-30,-20,49,-7,-55,46,40,-89,7,127,-113,-155,522,1023,522,-155,-113,127,7,-89,40,46,-55,-7,49,-20,-30,34,7,-34,12,23,-24,-7,26,-8,-19,18,7,-20,5,16,-14,-7,17,-3,-14,11,7,-14,2,12,-9,-7,12,-1,-11,7,6,-10,0,10,-6,-6,9,1,-9,5,6,-8,-1,8,-4,-6,7,2,-7,3,5,-6,-2,7,-2,-5,5,2,-6,2,5,-4,-2,5,-1,-5,4,2,-5,1,4,-3,-2,4,0,-4,3,2,-4,0,4,-2,-2,4,0,-4,2,2,-3,0,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm  Blackman-Harris de Nuttall 12
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-2,-1,2,0,-3,2,2,-3,0,3,-2,-2,3,0,-4,2,3,-3,-1,4,-2,-3,4,1,-5,2,4,-4,-2,5,-2,-5,4,2,-6,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-6,-5,9,0,-9,6,6,-10,-1,11,-6,-8,12,2,-13,6,10,-13,-3,16,-7,-13,15,5,-20,7,17,-18,-8,25,-7,-23,23,12,-33,7,34,-30,-20,49,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,49,-20,-30,34,7,-33,12,23,-23,-7,25,-8,-18,17,7,-20,5,15,-13,-7,16,-3,-13,10,6,-13,2,12,-8,-6,11,-1,-10,6,6,-9,0,9,-5,-6,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-6,2,4,-5,-2,5,-2,-4,4,2,-5,1,4,-3,-2,4,-1,-3,3,2,-4,0,3,-2,-2,3,0,-3,2,2,-3,0,2,-1,-2,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Parzen 13 
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,2,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,2,1,-2,0,2,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-4,2,3,-4,-1,4,-2,-3,4,1,-5,2,4,-4,-2,6,-2,-5,5,2,-6,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-6,-5,9,0,-10,6,7,-10,-1,11,-6,-8,12,2,-13,6,10,-13,-3,16,-7,-13,15,5,-20,7,17,-18,-8,25,-7,-23,23,12,-33,7,34,-30,-20,48,-7,-55,46,40,-88,7,127,-113,-155,522,1023,522,-155,-113,127,7,-88,40,46,-55,-7,48,-20,-30,34,7,-33,12,23,-23,-7,25,-8,-18,17,7,-20,5,15,-13,-7,16,-3,-13,10,6,-13,2,12,-8,-6,11,-1,-10,7,6,-10,0,9,-5,-6,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-6,2,5,-5,-2,6,-2,-4,4,2,-5,1,4,-3,-2,4,-1,-4,3,2,-4,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,2,0,-2,1,2,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,2,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Tukey 14
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-3,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,-1,-3,2,2,-3,0,3,-2,-2,4,0,-4,2,2,-4,0,4,-2,-3,4,0,-4,2,3,-4,-1,4,-2,-3,4,1,-5,2,4,-4,-1,5,-1,-4,4,2,-5,1,4,-4,-2,5,-1,-5,4,3,-5,0,5,-4,-3,6,0,-6,3,4,-6,0,6,-3,-4,6,1,-6,3,5,-6,-1,7,-3,-5,6,2,-7,3,6,-6,-3,8,-2,-7,6,3,-9,2,8,-7,-4,9,-1,-9,7,5,-10,1,10,-7,-6,11,0,-11,7,8,-12,-1,13,-7,-9,13,2,-15,7,12,-15,-3,18,-7,-14,16,5,-21,7,18,-19,-8,26,-7,-24,23,12,-34,7,34,-30,-20,49,-7,-55,46,40,-89,7,128,-113,-155,522,1023,522,-155,-113,128,7,-89,40,46,-55,-7,49,-20,-30,34,7,-34,12,23,-24,-7,26,-8,-19,18,7,-21,5,16,-14,-7,18,-3,-15,12,7,-15,2,13,-9,-7,13,-1,-12,8,7,-11,0,11,-6,-7,10,1,-10,5,7,-9,-1,9,-4,-7,8,2,-9,3,6,-7,-2,8,-3,-6,6,3,-7,2,6,-5,-3,7,-1,-6,5,3,-6,1,6,-4,-3,6,0,-6,4,3,-6,0,6,-3,-4,5,0,-5,3,4,-5,-1,5,-2,-4,4,1,-5,2,4,-4,-1,5,-1,-4,4,2,-5,1,4,-3,-2,4,-1,-4,3,2,-4,0,4,-3,-2,4,0,-4,2,2,-4,0,4,-2,-2,3,0,-3,2,2,-3,-1,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-3,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Triangular 15
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-4,2,2,-4,0,4,-2,-3,4,1,-4,2,3,-4,-1,5,-2,-4,4,1,-5,2,4,-5,-2,6,-2,-5,5,2,-7,1,6,-5,-3,7,-1,-7,5,4,-8,1,8,-5,-5,9,0,-9,6,6,-10,-1,11,-6,-8,11,2,-13,6,10,-13,-3,15,-6,-13,15,5,-19,7,17,-17,-7,24,-7,-22,22,12,-32,7,32,-29,-20,47,-7,-53,44,39,-87,7,126,-112,-153,520,1023,520,-153,-112,126,7,-87,39,44,-53,-7,47,-20,-29,32,7,-32,12,22,-22,-7,24,-7,-17,17,7,-19,5,15,-13,-6,15,-3,-13,10,6,-13,2,11,-8,-6,11,-1,-10,6,6,-9,0,9,-5,-5,8,1,-8,4,5,-7,-1,7,-3,-5,6,1,-7,2,5,-5,-2,6,-2,-5,4,2,-5,1,4,-4,-2,5,-1,-4,3,2,-4,1,4,-3,-2,4,0,-4,2,2,-4,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
		-- L=512 RANGE -1024 TO 1023 ofdm Retangular 16
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	-1,-2,2,1,-2,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,3,-1,-2,2,1,-2,1,2,-2,-1,3,-1,-2,2,1,-3,1,2,-2,-1,3,0,-2,2,1,-3,0,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-3,-1,4,0,-3,3,2,-4,0,4,-2,-2,4,0,-4,2,2,-4,0,4,-2,-3,4,1,-4,2,3,-4,-1,4,-2,-3,4,1,-4,2,4,-4,-1,5,-1,-4,4,2,-5,1,4,-4,-2,5,-1,-5,4,3,-5,1,5,-3,-3,6,0,-6,3,4,-6,0,6,-3,-4,6,1,-6,3,5,-6,-1,7,-3,-5,6,2,-7,3,6,-6,-2,8,-2,-7,7,3,-9,2,8,-7,-4,9,-1,-9,7,5,-10,1,10,-7,-6,11,0,-11,7,8,-12,-1,13,-7,-9,13,2,-15,7,12,-14,-3,18,-7,-14,17,5,-21,7,18,-19,-8,26,-7,-24,23,13,-34,7,34,-30,-20,49,-7,-55,46,40,-89,7,128,-113,-155,522,1023,522,-155,-113,128,7,-89,40,46,-55,-7,49,-20,-30,34,7,-34,13,23,-24,-7,26,-8,-19,18,7,-21,5,17,-14,-7,18,-3,-14,12,7,-15,2,13,-9,-7,13,-1,-12,8,7,-11,0,11,-6,-7,10,1,-10,5,7,-9,-1,9,-4,-7,8,2,-9,3,7,-7,-2,8,-2,-6,6,3,-7,2,6,-5,-3,7,-1,-6,5,3,-6,1,6,-4,-3,6,0,-6,4,3,-6,0,6,-3,-3,5,1,-5,3,4,-5,-1,5,-2,-4,4,1,-5,2,4,-4,-1,5,-1,-4,4,2,-4,1,4,-3,-2,4,-1,-4,3,2,-4,1,4,-3,-2,4,0,-4,2,2,-4,0,4,-2,-2,4,0,-4,2,3,-3,0,4,-1,-3,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,3,0,-3,1,2,-2,0,3,-1,-2,2,1,-3,1,2,-2,-1,3,-1,-2,2,1,-2,1,2,-2,-1,3,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,0,2,-1,-2,2,1,-2,1,2,-2,-1,2
	--);
	-- >>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>

	-- L=1024 RANGE -512 TO 511 ofdm hamming
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,0,0,0,0,1,0,0,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,-1,2,-1,-2,2,1,-2,0,2,-2,-1,2,0,-2,2,1,-2,0,2,-2,-1,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,1,2,-3,-1,3,-1,-3,3,1,-4,1,3,-3,-1,4,-1,-3,3,2,-4,1,4,-3,-2,5,-1,-4,3,2,-5,0,5,-3,-3,5,0,-6,3,4,-6,0,6,-3,-5,6,1,-7,4,6,-7,-2,9,-4,-7,8,3,-10,4,9,-10,-4,13,-4,-12,12,6,-17,4,17,-15,-10,24,-4,-27,23,20,-44,4,64,-56,-77,261,511,261,-77,-56,64,4,-44,20,23,-27,-4,24,-10,-15,17,4,-17,6,12,-12,-4,13,-4,-10,9,4,-10,3,8,-7,-4,9,-2,-7,6,4,-7,1,6,-5,-3,6,0,-6,4,3,-6,0,5,-3,-3,5,0,-5,2,3,-4,-1,5,-2,-3,4,1,-4,2,3,-3,-1,4,-1,-3,3,1,-4,1,3,-3,-1,3,-1,-3,2,1,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-1,-2,2,0,-2,1,2,-2,0,2,-1,-2,2,0,-2,1,2,-2,-1,2,-1,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,0,0,1,0,0,0,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=2048 RANGE -127 to 126 HAMMING
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,4,4,4,4,4,4,4,3,3,3,3,3,3,2,2,2,2,2,1,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-3,-4,-4,-4,-4,-5,-5,-5,-5,-5,-6,-6,-6,-6,-6,-7,-7,-7,-7,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-8,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-8,-8,-8,-8,-8,-8,-8,-8,-7,-7,-7,-7,-7,-6,-6,-6,-6,-5,-5,-5,-5,-4,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,0,0,0,1,1,1,2,2,2,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,11,12,12,12,12,12,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,13,13,13,13,13,12,12,12,12,11,11,11,10,10,10,9,9,9,8,8,7,7,6,6,5,5,4,4,3,3,2,2,1,1,0,-1,-1,-2,-2,-3,-4,-4,-5,-6,-6,-7,-7,-8,-9,-9,-10,-11,-11,-12,-12,-13,-14,-14,-15,-15,-16,-16,-17,-18,-18,-19,-19,-20,-20,-21,-21,-22,-22,-22,-23,-23,-24,-24,-24,-25,-25,-25,-25,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-25,-25,-25,-25,-24,-24,-24,-23,-23,-22,-22,-21,-21,-20,-19,-19,-18,-17,-16,-16,-15,-14,-13,-12,-11,-10,-9,-8,-7,-6,-5,-4,-2,-1,0,1,2,4,5,6,8,9,11,12,14,15,17,18,20,21,23,24,26,28,29,31,33,34,36,38,39,41,43,44,46,48,50,51,53,55,57,58,60,62,64,65,67,69,70,72,74,75,77,79,80,82,84,85,87,88,90,91,93,94,96,97,99,100,101,103,104,105,106,108,109,110,111,112,113,114,115,116,117,118,119,120,120,121,122,122,123,123,124,124,125,125,126,126,126,126,127,127,127,127,127,127,127,127,126,126,126,126,125,125,124,124,123,123,122,122,121,120,120,119,118,117,116,115,114,113,112,111,110,109,108,106,105,104,103,101,100,99,97,96,94,93,91,90,88,87,85,84,82,80,79,77,75,74,72,70,69,67,65,64,62,60,58,57,55,53,51,50,48,46,44,43,41,39,38,36,34,33,31,29,28,26,24,23,21,20,18,17,15,14,12,11,9,8,6,5,4,2,1,0,-1,-2,-4,-5,-6,-7,-8,-9,-10,-11,-12,-13,-14,-15,-16,-16,-17,-18,-19,-19,-20,-21,-21,-22,-22,-23,-23,-24,-24,-24,-25,-25,-25,-25,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-25,-25,-25,-25,-24,-24,-24,-23,-23,-22,-22,-22,-21,-21,-20,-20,-19,-19,-18,-18,-17,-16,-16,-15,-15,-14,-14,-13,-12,-12,-11,-11,-10,-9,-9,-8,-7,-7,-6,-6,-5,-4,-4,-3,-2,-2,-1,-1,0,1,1,2,2,3,3,4,4,5,5,6,6,7,7,8,8,9,9,9,10,10,10,11,11,11,12,12,12,12,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,13,13,13,13,13,12,12,12,12,12,11,11,11,11,10,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,2,2,2,1,1,1,0,0,0,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-4,-5,-5,-5,-5,-6,-6,-6,-6,-7,-7,-7,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-8,-8,-8,-8,-8,-8,-8,-8,-8,-7,-7,-7,-7,-7,-7,-6,-6,-6,-6,-6,-5,-5,-5,-5,-5,-4,-4,-4,-4,-3,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,1,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,3,3,3,3,3,3,3,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- degrau tamanho 512
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	0,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- rect tamanho 512, valor 100 do índice 56 até o 512-56 (pulso de tamanho 400)
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- degrau tamanho 1024
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	0,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- noisy sin -127 to 126
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-10,1,11,35,36,18,49,41,42,51,51,56,70,75,79,79,72,87,96,93,100,
	--	101,98,104,100,111,101,103,106,95,121,115,109,121,103,111,109,111,
	--	110,101,104,101,103,103,100,85,87,76,73,75,80,62,64,56,59,41,42,40,
	--	38,35,21,6,5,-3,11,-11,-9,-20,-19,-35,-44,-49,-43,-52,-58,-53,-64,
	--	-70,-66,-84,-80,-83,-93,-93,-105,-108,-103,-102,-94,-114,-111,-114,
	--	-126,-119,-127,-112,-122,-117,-120,-114);

	--noisy sawtooth -64 to 63
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-30,-25,-33,-32,-20,-46,-30,-35,-26,-15,-12,-27,-20,-13,-15,-8 ,-6 ,-16,-8 ,-24,7  ,-7 ,-11,0  ,-9 ,5  ,2  ,28 ,20 ,-11,17 ,2  ,14 ,19 ,26 ,19 ,37 ,20 ,29 ,33 ,30 ,39 ,35 ,27 ,19 ,54 ,33 ,41 ,47 ,44 ,37 ,42 ,47 ,63 ,44 ,60 ,57 ,54 ,48 ,57 ,60 ,50 ,-35,-42,-34,-29,-38,-31,-24,-42,-14,0  ,-12,-22,-13,-25,3  ,-4 ,-4 ,-17,-5 ,-11,-7 ,-8 ,-10,-8 ,0  ,-12,11 ,6  ,15 ,13 ,16 ,0  ,6  ,12 ,19 ,30 ,19 ,34
	--	);

	--noisy sawtooth -256 to 255
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-155,-124,-155,-177,-200,-134,-104,-138,-140,-125,-147,-119,-102,-87 ,-85 ,-54 ,-65 ,2   ,-45 ,15  ,-70 ,-18 ,-40 ,-3  ,3   ,-90 ,-53 ,-50 ,22  ,67  ,9   ,56  ,53  ,2   ,61  ,26  ,114 ,64  ,131 ,63  ,106 ,89  ,25  ,69  ,133 ,115 ,83  ,107 ,145 ,107 ,184 ,132 ,227 ,130 ,182 ,127 ,162 ,173 ,215 ,241 ,224 ,206 ,256 ,-142,-160,-138,-137,-181,-112,-156,-148,-113,-124,-112,-79 ,-56 ,-95 ,-69 ,-83 ,-60 ,-46 ,-78 ,-39 ,-21 ,-33 ,32  ,-45 ,-43 ,-73 ,29  ,34  ,6   ,48  ,28  ,39  ,39  ,57  ,51  ,154 ,18		
	--);

	-- TAMANHO 1060 - Símbolo OFDM parte real, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,-8,-252,-50,257,131,-90,5,157,127,28,-93,-149,13,112,-163,-382,-122,189,158,75,50,-166,-386,-280,-62,56,178,156,-138,-239,35,83,-201,-143,231,201,-134,-148,1,-117,-248,-126,-9,2,87,129,-59,-271,-297,-202,-33,141,83,-163,-215,-66,-97,-263,-163,123,159,-20,-31,131,200,217,341,368,100,-137,-28,131,38,-18,179,270,60,-114,-110,-115,-81,52,-8,-247,-187,132,176,39,121,92,-338,-512,-44,336,189,63,176,112,-90,-67,20,-13,69,172,-87,-376,-133,229,58,-304,-288,-133,-161,-152,-17,-24,-148,-149,-103,-160,-203,-158,-129,-90,43,175,221,202,51,-220,-289,-14,210,91,-72,3,85,-48,-167,-25,196,187,-7,-75,77,226,197,58,-77,-135,-26,191,227,19,-99,13,48,-119,-185,-14,138,105,-7,-104,-172,-151,2,184,210,29,-159,-169,-116,-120,-8,225,186,-104,-43,339,272,-225,-285,114,187,-14,158,477,337,16,45,179,45,-156,-171,-75,31,77,-34,-202,-229,-164,-112,-2,112,34,-119,-49,160,181,4,-106,-8,186,250,115,-8,-1,-61,-202,-102,179,155,-121,-81,239,290,115,159,267,41,-228,-63,287,284,-20,-204,-157,-101,-174,-232,-56,255,328,94,-53,36,11,-217,-228,49,140,-45,-60,109,12,-313,-394,-226,-153,-178,-138,-96,-73,16,11,-215,-365,-244,-130,-145,-76,-21,-204,-296,-6,207,-5,-209,-135,-115,-189,-86,-34,-244,-209,268,447,71,-90,178,183,-131,-134,82,-16,-223,-157,-133,-348,-375,-130,-45,-77,99,201,-86,-292,-7,338,313,117,-46,-220,-281,-96,99,58,-109,-215,-183,-6,125,-24,-241,-108,242,305,42,-131,-13,202,265,149,52,97,127,35,-9,56,57,36,179,300,140,-77,-95,-73,-87,46,211,125,-25,51,150,39,-51,65,170,68,-127,-204,-96,53,96,145,303,322,100,17,194,195,-36,-18,230,190,-114,-226,-86,105,261,236,-21,-195,-152,-181,-259,-17,368,361,41,-120,-67,-9,-6,-78,-192,-174,-20,54,55,143,232,174,56,-12,-31,-25,-94,-263,-259,57,301,220,109,115,43,-34,58,80,-61,3,278,314,123,46,8,-77,3,84,-165,-312,105,468,163,-240,-149,16,-107,-151,49,138,24,-13,76,92,-11,-104,-147,-217,-276,-153,82,98,-75,-58,66,-105,-355,-225,-21,-172,-298,-93,-26,-247,-185,209,309,60,-46,9,-52,-124,-38,49,49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- TAMANHO 1060 - Símbolo OFDM parte imaginária, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,-241,-142,-79,-110,-46,-71,-296,-384,-232,-109,17,300,443,217,-3,66,131,-16,-132,-64,31,78,150,181,59,-55,59,201,8,-327,-267,80,90,-225,-240,70,115,-147,-184,64,136,-73,-201,-68,116,121,0,-46,19,12,-155,-341,-401,-342,-250,-197,-172,-110,-78,-175,-203,51,280,108,-189,-172,11,80,137,199,80,-51,88,265,191,87,129,79,-124,-203,-104,-26,-33,-85,-129,-47,129,164,58,44,92,53,53,139,59,-177,-251,-176,-158,-81,88,14,-268,-254,66,195,108,138,211,138,91,111,-100,-466,-465,-32,262,78,-250,-268,-3,153,26,-161,-198,-138,-45,63,35,-146,-126,222,407,129,-168,-117,-36,-211,-380,-298,-89,106,239,191,-11,-91,29,102,24,-58,-112,-179,-112,128,206,-49,-245,-59,190,133,-14,73,212,114,-108,-231,-248,-160,38,128,-31,-134,26,87,-180,-350,-147,-1,-217,-432,-339,-134,-5,125,246,217,47,-112,-151,-115,-150,-249,-210,-77,-146,-270,1,405,262,-189,-178,118,30,-220,-79,180,106,-79,-106,-112,-141,-93,-51,-13,198,425,308,-20,-125,29,162,122,-38,-135,-34,128,186,215,202,4,-107,199,465,137,-321,-258,49,127,67,-36,-198,-147,139,143,-155,-187,-4,-83,-227,-121,-98,-266,-193,34,-35,-163,6,139,66,144,279,76,-185,-129,-73,-194,-162,-40,-181,-347,-180,102,270,382,335,142,165,312,96,-219,-43,238,11,-296,-145,99,97,97,106,-101,-281,-154,1,-66,-142,-47,142,258,89,-318,-436,-27,333,196,-58,-33,86,98,61,-7,-83,-31,102,105,-3,-60,-55,-31,-10,-72,-175,-106,94,120,-28,-69,-15,-49,-51,124,265,197,122,168,114,-152,-357,-266,-73,-69,-142,35,376,419,67,-220,-125,122,213,154,76,51,108,171,117,12,36,128,87,-17,32,175,182,32,-132,-231,-230,-128,-16,67,138,56,-250,-368,3,302,-23,-363,13,511,294,-139,22,371,226,-92,-65,70,9,-45,59,143,127,98,97,136,167,34,-227,-286,-46,137,26,-140,-81,110,140,-56,-232,-165,50,170,133,23,-87,-110,-14,66,45,69,205,223,-28,-320,-322,2,349,374,100,-83,5,79,-58,-176,-73,124,234,216,98,-15,-33,-59,-171,-187,-22,53,-71,-95,90,156,-9,-79,48,69,-82,-88,92,94,-162,-316,-222,-113,-105,-108,-92,-7,200,271,-5,-199,70,278,-47,-332,-62,265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- A saída da convolução vai ter tamanho 1572

	-- TAMANHO 1060 - Símbolo OFDM parte real, -1024 to 1023
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	97,213,470,554,368,99,-75,-138,-167,-126,10,-63,-548,-931,-650,-34,246,143,34,99,196,68,-202,-139,221,205,-161,-76,428,620,556,552,211,-348,-240,237,-17,-504,-99,513,263,-180,10,314,253,56,-186,-298,26,225,-325,-764,-243,378,316,150,100,-333,-771,-561,-123,113,356,311,-275,-478,69,166,-403,-285,463,402,-269,-295,2,-234,-497,-251,-17,3,174,258,-118,-543,-594,-404,-65,282,166,-326,-430,-131,-194,-527,-326,246,318,-41,-63,262,400,434,682,735,201,-274,-56,263,76,-36,358,539,120,-228,-220,-230,-162,103,-15,-495,-373,265,352,78,242,185,-676,-1024,-88,671,379,126,352,224,-179,-135,40,-27,138,344,-174,-751,-266,458,115,-607,-576,-266,-323,-303,-34,-47,-295,-299,-207,-321,-405,-315,-257,-180,85,350,442,404,102,-439,-578,-28,421,183,-144,5,170,-96,-333,-50,392,373,-13,-150,154,452,394,115,-153,-271,-51,383,455,38,-198,25,96,-237,-370,-29,276,210,-14,-207,-343,-302,3,368,419,59,-317,-339,-232,-241,-16,450,371,-208,-86,678,543,-451,-571,228,374,-28,316,955,673,32,90,359,90,-313,-343,-151,62,154,-68,-403,-458,-328,-224,-4,224,68,-238,-97,320,362,9,-211,-16,373,500,229,-15,-1,-121,-403,-204,358,309,-241,-162,479,581,230,319,534,83,-456,-125,574,569,-39,-408,-315,-202,-348,-464,-112,511,655,188,-107,72,22,-434,-457,99,279,-91,-121,219,23,-627,-789,-451,-306,-356,-275,-193,-146,32,22,-431,-731,-487,-260,-290,-152,-43,-409,-593,-13,414,-10,-418,-271,-231,-378,-173,-68,-489,-418,536,894,142,-181,356,366,-262,-268,164,-33,-446,-314,-266,-697,-750,-260,-90,-154,199,402,-172,-584,-14,676,627,233,-92,-440,-563,-192,197,116,-219,-430,-366,-13,250,-48,-482,-216,483,609,83,-262,-25,405,530,298,105,194,254,71,-18,112,114,73,359,599,280,-155,-190,-146,-174,93,421,250,-50,103,299,77,-102,131,340,136,-254,-408,-193,105,191,291,605,645,201,34,388,390,-73,-36,459,380,-227,-452,-172,211,523,472,-42,-391,-305,-362,-518,-34,736,722,82,-240,-133,-19,-13,-155,-384,-347,-40,109,110,285,464,349,111,-24,-61,-50,-187,-527,-517,115,602,441,217,231,87,-67,115,160,-123,6,557,628,247,92,16,-154,6,167,-329,-623,210,936,325,-480,-299,32,-213,-302,98,275,47,-26,152,184,-21,-207,-293,-433,-552,-305,165,197,-150,-117,133,-210,-709,-450,-42,-343,-595,-186,-52,-495,-370,419,619,120,-92,19,-105,-248,-76,97,97,213,470,554,368,99,-75,-138,-167,-126,10,-63,-548,-931,-650,-34,246,143,34,99,196,68,-202,-139,221,205,-161,-76,428,620,556,552,211,-348,-240,237,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- TAMANHO 1060 - Símbolo OFDM parte imaginária, -1024 to 1023
	constant NOISY_ARRAY : T_NOISY_INPUT := (
		530,470,334,262,-238,-476,236,783,330,-60,175,119,-249,17,584,518,136,4,-97,-103,275,438,-82,-500,-239,111,103,-27,-101,-3,282,221,-319,-358,399,681,0,-482,-285,-158,-221,-92,-142,-592,-768,-465,-218,35,601,886,434,-7,131,262,-31,-264,-128,62,155,300,362,118,-109,118,403,16,-654,-536,159,179,-450,-480,141,230,-295,-369,128,272,-146,-403,-136,231,243,0,-91,38,24,-311,-682,-802,-685,-500,-394,-344,-220,-156,-350,-406,102,561,216,-379,-344,21,159,274,398,160,-102,175,530,383,173,258,159,-248,-406,-208,-52,-67,-170,-258,-94,258,328,117,88,184,106,106,278,118,-355,-502,-352,-317,-163,177,29,-537,-508,132,391,217,276,422,276,181,222,-200,-933,-931,-63,525,156,-501,-536,-7,306,51,-322,-397,-277,-90,127,70,-293,-253,444,815,258,-337,-234,-72,-423,-761,-596,-179,212,478,381,-22,-182,59,205,48,-117,-225,-358,-224,255,412,-99,-490,-118,381,265,-27,146,425,229,-216,-463,-497,-321,77,256,-62,-268,51,174,-361,-700,-294,-2,-434,-866,-678,-269,-11,251,492,434,94,-223,-302,-230,-300,-498,-421,-155,-292,-541,3,812,525,-378,-356,236,59,-440,-158,360,213,-159,-212,-223,-283,-187,-102,-26,397,851,616,-40,-250,59,325,245,-77,-271,-68,257,372,430,404,8,-214,399,930,275,-642,-517,98,254,133,-71,-397,-293,278,286,-310,-374,-9,-166,-454,-242,-196,-533,-387,67,-71,-326,12,279,131,288,558,151,-370,-259,-145,-389,-324,-80,-361,-694,-360,205,541,765,670,284,331,626,193,-439,-86,476,21,-593,-290,197,195,194,213,-202,-563,-308,1,-132,-284,-93,284,517,177,-637,-873,-54,667,393,-115,-67,173,196,122,-13,-165,-62,203,211,-6,-121,-110,-62,-20,-143,-350,-212,188,240,-56,-139,-30,-98,-102,249,530,395,244,336,229,-305,-714,-532,-146,-138,-284,70,752,839,133,-439,-250,244,427,309,152,102,216,342,234,24,72,256,175,-33,65,350,364,65,-264,-463,-461,-257,-31,134,277,112,-500,-738,6,605,-46,-727,25,1023,588,-278,43,743,452,-184,-131,139,17,-89,118,287,254,196,195,273,335,68,-455,-573,-93,273,52,-281,-161,219,280,-112,-464,-329,99,339,266,45,-174,-220,-28,133,90,137,409,447,-56,-640,-645,3,699,748,199,-165,11,157,-116,-353,-146,248,469,433,196,-30,-66,-118,-343,-373,-44,106,-143,-191,179,312,-17,-159,96,138,-164,-175,185,188,-324,-633,-445,-226,-210,-216,-185,-14,401,543,-11,-399,139,557,-93,-665,-125,530,470,334,262,-238,-476,236,783,330,-60,175,119,-249,17,584,518,136,4,-97,-103,275,438,-82,-500,-239,111,103,-27,-101,-3,282,221,-319,-358,399,681,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);
	-- A saída da convolução vai ter tamanho 1572

	-- TAMANHO 1572 - Símbolo OFDM parte real, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,-8,-252,-50,257,131,-90,5,157,127,28,-93,-149,13,112,-163,-382,-122,189,158,75,50,-166,-386,-280,-62,56,178,156,-138,-239,35,83,-201,-143,231,201,-134,-148,1,-117,-248,-126,-9,2,87,129,-59,-271,-297,-202,-33,141,83,-163,-215,-66,-97,-263,-163,123,159,-20,-31,131,200,217,341,368,100,-137,-28,131,38,-18,179,270,60,-114,-110,-115,-81,52,-8,-247,-187,132,176,39,121,92,-338,-512,-44,336,189,63,176,112,-90,-67,20,-13,69,172,-87,-376,-133,229,58,-304,-288,-133,-161,-152,-17,-24,-148,-149,-103,-160,-203,-158,-129,-90,43,175,221,202,51,-220,-289,-14,210,91,-72,3,85,-48,-167,-25,196,187,-7,-75,77,226,197,58,-77,-135,-26,191,227,19,-99,13,48,-119,-185,-14,138,105,-7,-104,-172,-151,2,184,210,29,-159,-169,-116,-120,-8,225,186,-104,-43,339,272,-225,-285,114,187,-14,158,477,337,16,45,179,45,-156,-171,-75,31,77,-34,-202,-229,-164,-112,-2,112,34,-119,-49,160,181,4,-106,-8,186,250,115,-8,-1,-61,-202,-102,179,155,-121,-81,239,290,115,159,267,41,-228,-63,287,284,-20,-204,-157,-101,-174,-232,-56,255,328,94,-53,36,11,-217,-228,49,140,-45,-60,109,12,-313,-394,-226,-153,-178,-138,-96,-73,16,11,-215,-365,-244,-130,-145,-76,-21,-204,-296,-6,207,-5,-209,-135,-115,-189,-86,-34,-244,-209,268,447,71,-90,178,183,-131,-134,82,-16,-223,-157,-133,-348,-375,-130,-45,-77,99,201,-86,-292,-7,338,313,117,-46,-220,-281,-96,99,58,-109,-215,-183,-6,125,-24,-241,-108,242,305,42,-131,-13,202,265,149,52,97,127,35,-9,56,57,36,179,300,140,-77,-95,-73,-87,46,211,125,-25,51,150,39,-51,65,170,68,-127,-204,-96,53,96,145,303,322,100,17,194,195,-36,-18,230,190,-114,-226,-86,105,261,236,-21,-195,-152,-181,-259,-17,368,361,41,-120,-67,-9,-6,-78,-192,-174,-20,54,55,143,232,174,56,-12,-31,-25,-94,-263,-259,57,301,220,109,115,43,-34,58,80,-61,3,278,314,123,46,8,-77,3,84,-165,-312,105,468,163,-240,-149,16,-107,-151,49,138,24,-13,76,92,-11,-104,-147,-217,-276,-153,82,98,-75,-58,66,-105,-355,-225,-21,-172,-298,-93,-26,-247,-185,209,309,60,-46,9,-52,-124,-38,49,49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- TAMANHO 1572 - Símbolo OFDM parte imaginária, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,-241,-142,-79,-110,-46,-71,-296,-384,-232,-109,17,300,443,217,-3,66,131,-16,-132,-64,31,78,150,181,59,-55,59,201,8,-327,-267,80,90,-225,-240,70,115,-147,-184,64,136,-73,-201,-68,116,121,0,-46,19,12,-155,-341,-401,-342,-250,-197,-172,-110,-78,-175,-203,51,280,108,-189,-172,11,80,137,199,80,-51,88,265,191,87,129,79,-124,-203,-104,-26,-33,-85,-129,-47,129,164,58,44,92,53,53,139,59,-177,-251,-176,-158,-81,88,14,-268,-254,66,195,108,138,211,138,91,111,-100,-466,-465,-32,262,78,-250,-268,-3,153,26,-161,-198,-138,-45,63,35,-146,-126,222,407,129,-168,-117,-36,-211,-380,-298,-89,106,239,191,-11,-91,29,102,24,-58,-112,-179,-112,128,206,-49,-245,-59,190,133,-14,73,212,114,-108,-231,-248,-160,38,128,-31,-134,26,87,-180,-350,-147,-1,-217,-432,-339,-134,-5,125,246,217,47,-112,-151,-115,-150,-249,-210,-77,-146,-270,1,405,262,-189,-178,118,30,-220,-79,180,106,-79,-106,-112,-141,-93,-51,-13,198,425,308,-20,-125,29,162,122,-38,-135,-34,128,186,215,202,4,-107,199,465,137,-321,-258,49,127,67,-36,-198,-147,139,143,-155,-187,-4,-83,-227,-121,-98,-266,-193,34,-35,-163,6,139,66,144,279,76,-185,-129,-73,-194,-162,-40,-181,-347,-180,102,270,382,335,142,165,312,96,-219,-43,238,11,-296,-145,99,97,97,106,-101,-281,-154,1,-66,-142,-47,142,258,89,-318,-436,-27,333,196,-58,-33,86,98,61,-7,-83,-31,102,105,-3,-60,-55,-31,-10,-72,-175,-106,94,120,-28,-69,-15,-49,-51,124,265,197,122,168,114,-152,-357,-266,-73,-69,-142,35,376,419,67,-220,-125,122,213,154,76,51,108,171,117,12,36,128,87,-17,32,175,182,32,-132,-231,-230,-128,-16,67,138,56,-250,-368,3,302,-23,-363,13,511,294,-139,22,371,226,-92,-65,70,9,-45,59,143,127,98,97,136,167,34,-227,-286,-46,137,26,-140,-81,110,140,-56,-232,-165,50,170,133,23,-87,-110,-14,66,45,69,205,223,-28,-320,-322,2,349,374,100,-83,5,79,-58,-176,-73,124,234,216,98,-15,-33,-59,-171,-187,-22,53,-71,-95,90,156,-9,-79,48,69,-82,-88,92,94,-162,-316,-222,-113,-105,-108,-92,-7,200,271,-5,-199,70,278,-47,-332,-62,265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- A saída da convolução vai ter tamanho 2596

-- in=2000, out=2000, seno + ruído aleatório (white gaussian noise) (converge mais ou menos)
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	-2,9,9,2,20,34,51,57,40,43,45,36,71,62,46,59,59,59,38,55,75,75,65,67,66,71,59,64,63,48,50,80,67,67,62,45,74,57,43,50,24,35,26,30,36,11,32,15,6,-1,5,-4,-12,-28,-28,-26,8,-22,-30,-42,-63,-40,-51,-38,-55,-71,-52,-66,-60,-60,-30,-68,-62,-71,-76,-73,-68,-58,-63,-56,-49,-54,-54,-60,-53,-36,-48,-40,-54,-12,-20,-34,-22,-20,-16,-19,8,-7,14,-15,22,-5,13,14,30,37,48,35,36,44,32,45,49,64,56,58,57,76,59,59,67,63,80,91,71,78,76,66,66,51,75,79,51,41,61,36,52,40,40,53,41,17,32,39,20,-4,27,8,2,20,1,-22,-14,-23,-26,-25,-40,-16,-39,-18,-23,-46,-56,-57,-51,-61,-59,-54,-70,-57,-36,-50,-66,-69,-57,-49,-46,-76,-45,-38,-66,-54,-63,-60,-39,-46,-45,-50,-55,-32,-27,-8,-32,-13,-16,3,-12,-17,6,-15,-2,27,21,28,48,23,36,28,51,35,61,47,39,37,57,39,46,63,72,73,58,66,42,53,79,73,69,45,63,75,70,59,56,61,73,40,61,51,28,26,45,17,25,42,31,5,25,4,12,2,17,-19,-28,-12,-2,-21,-23,-13,-41,-48,-34,-29,-53,-13,-51,-68,-55,-64,-81,-58,-82,-58,-25,-66,-84,-62,-64,-64,-66,-73,-65,-80,-83,-50,-43,-31,-52,-24,-22,-27,-34,-23,-39,-37,-40,-8,-15,-4,10,-1,1,15,24,27,25,13,23,13,44,46,60,44,60,52,45,45,68,73,56,56,67,71,85,85,70,68,74,71,50,58,69,54,50,50,57,67,49,37,57,31,24,41,19,26,44,23,12,21,-16,2,-0,3,2,-8,-26,-14,-22,-37,-24,-48,-30,-37,-52,-47,-59,-65,-36,-58,-46,-45,-68,-65,-52,-48,-72,-67,-82,-78,-72,-70,-58,-53,-43,-36,-37,-59,-31,-30,-58,-37,-8,-40,-28,-25,-20,-6,-0,-2,-8,10,-11,15,12,7,33,27,36,7,57,44,8,51,36,48,59,73,80,64,55,72,54,57,56,59,74,57,72,73,48,72,52,61,54,55,55,48,42,65,62,45,34,22,24,15,28,2,22,20,3,5,-17,-13,-3,-26,-11,-22,-15,-29,-23,-51,-37,-24,-52,-38,-50,-40,-67,-65,-68,-35,-70,-71,-51,-70,-73,-60,-44,-98,-47,-44,-12,-51,-63,-62,-47,-42,-54,-56,-47,-31,-35,-16,-25,-32,-15,-26,-20,16,-4,11,3,-5,-2,25,21,5,35,50,46,44,62,50,61,66,48,66,67,57,76,58,63,75,72,82,51,45,70,56,69,75,50,53,61,26,67,52,69,48,33,32,48,20,40,25,26,30,34,5,-3,19,-2,2,-20,-17,-31,-23,-30,-15,-37,-23,-46,-59,-52,-53,-65,-71,-38,-49,-57,-48,-82,-57,-70,-63,-60,-61,-56,-74,-63,-68,-47,-66,-63,-51,-66,-30,-49,-47,-43,-37,-13,-33,-40,-7,-20,-24,-27,-7,14,-1,8,-6,-9,18,32,6,32,47,53,34,69,35,48,51,72,48,48,55,61,90,67,66,70,71,71,68,46,82,42,68,64,59,67,77,54,69,55,59,42,29,38,33,28,20,33,25,26,36,-1,-6,10,1,-4,-4,-21,-3,-30,-36,-19,-48,-24,-41,-33,-48,-26,-68,-51,-58,-58,-60,-58,-56,-66,-60,-51,-60,-55,-61,-36,-62,-64,-70,-61,-52,-54,-39,-37,-29,-58,-19,-36,-16,-14,-13,-6,-20,-16,-7,12,-1,-6,9,17,14,18,37,35,34,39,42,46,50,37,89,43,77,47,57,69,31,43,58,75,62,71,63,61,63,74,68,62,76,66,60,52,54,51,51,37,36,25,32,5,34,43,-3,23,-3,19,-22,-12,10,-3,-3,-18,-21,-37,-11,-32,-34,-7,-53,-52,-43,-32,-50,-40,-62,-51,-40,-77,-69,-70,-78,-72,-77,-67,-47,-46,-59,-71,-63,-41,-59,-36,-30,-57,-45,-36,-39,-35,1,-51,-11,-22,-18,-12,29,-15,9,14,-9,1,24,20,19,9,45,17,44,48,67,58,60,67,80,74,54,57,67,100,54,57,55,57,66,76,71,57,60,51,53,63,60,68,68,34,35,40,35,30,32,22,32,15,13,4,21,6,-6,6,-4,-23,5,-22,-22,-7,-21,-33,-27,-51,-38,-45,-57,-52,-55,-26,-87,-67,-36,-50,-61,-62,-55,-67,-60,-80,-49,-65,-54,-64,-27,-70,-35,-20,-54,-27,-57,-41,-21,-43,-38,-29,-26,-31,-19,-14,-14,9,-18,20,23,25,-2,40,21,28,38,50,51,48,53,52,38,60,78,45,62,54,70,71,58,65,65,57,52,44,65,71,81,56,65,67,63,64,64,62,53,38,36,46,45,23,16,21,26,7,20,-10,33,3,-24,-12,-21,-29,-40,-38,-22,-27,-20,-36,-48,-62,-34,-53,-72,-40,-60,-54,-63,-80,-37,-88,-68,-67,-61,-76,-53,-50,-59,-94,-59,-50,-51,-72,-38,-49,-32,-39,-30,-19,-20,-18,-25,4,-32,-4,-7,-7,-8,9,25,23,15,30,26,17,25,17,46,54,32,36,64,59,44,58,76,88,68,49,72,64,83,70,58,69,63,92,49,55,52,56,64,58,56,72,64,46,25,37,24,10,37,32,30,10,-10,-15,-12,-6,8,-12,-3,-21,-23,-12,-38,-32,-28,-59,-45,-42,-31,-51,-46,-49,-73,-68,-48,-48,-61,-64,-66,-48,-71,-64,-77,-59,-49,-58,-63,-54,-63,-32,-56,-26,-36,-29,-21,-39,-33,-20,-38,-21,8,-20,-13,6,1,19,16,12,25,38,23,39,31,37,58,38,62,59,65,75,45,72,60,47,99,67,67,81,72,57,34,69,71,68,62,61,75,53,67,40,46,56,47,52,41,43,31,24,18,15,-5,-2,-7,-6,21,-21,-25,-17,-13,2,-29,-40,-28,-31,-34,-30,-56,-38,-63,-40,-69,-61,-52,-74,-60,-58,-58,-46,-88,-66,-53,-94,-53,-49,-69,-61,-58,-54,-41,-58,-30,-59,-51,-36,-33,-34,-20,-29,-39,-32,-7,-25,-26,9,-10,2,29,11,42,24,1,25,49,50,31,27,53,35,58,54,64,50,67,68,81,75,59,73,84,71,51,77,75,58,85,67,71,49,69,25,63,61,56,43,49,29,9,41,26,12,15,19,10,7,9,6,-24,-37,-18,-16,-17,-13,-24,-38,-54,-36,-53,-45,-44,-35,-39,-44,-45,-57,-57,-74,-40,-70,-59,-46,-64,-51,-61,-58,-56,-69,-75,-59,-35,-39,-40,-53,-33,-19,-60,-42,-26,-19,-1,-34,-1,1,6,6,24,12,-15,16,33,14,34,28,27,33,33,42,51,56,68,62,63,54,65,71,49,70,58,82,74,82,68,86,72,72,58,55,82,60,60,52,31,45,36,38,49,46,39,29,29,43,18,18,2,9,-21,4,8,2,-36,-27,-11,-23,-19,-41,-29,-43,-35,-33,-47,-46,-43,-68,-58,-43,-49,-71,-65,-59,-49,-68,-75,-60,-64,-67,-65,-58,-69,-90,-50,-34,-24,-65,-47,-48,-16,-38,-34,-17,-3,-14,-1,-15,-21,-9,8,-2,19,30,21,33,38,22,39,48,40,41,69,52,56,79,46,50,44,50,76,40,76,76,70,44,77,83,75,62,65,68,93,66,72,43,55,40,54,24,32,26,32,59,21,40,14,32,-9,-3,7,8,3,-10,-25,-16,-19,-37,-19,-36,-11,-23,-32,-53,-75,-47,-60,-41,-41,-82,-65,-55,-66,-84,-42,-56,-56,-71,-46,-45,-61,-73,-60,-50,-59,-62,-22,-42,-36,-57,-34,-24,-42,-14,-5,-15,-8,-13,-5,-3,16,17,14,10,42,41,33,40,27,45,40,50,62,58,57,53,57,65,59,64,65,72,48,94,76,57,75,44,55,69,72,65,78,63,49,41,45,42,56,57,33,44,46,52,44,3,23,31,-7,9,16,1,-18,-14,-14,-12,-13,-40,-10,-49,-33,-34,-25,-52,-36,-69,-58,-41,-46,-49,-59,-55,-67,-58,-82,-68,-62,-56,-100,-57,-69,-68,-34,-58,-39,-47,-42,-46,-51,-57,-32,-36,-53,-30,-44,-16,-6,-17,-1,17,9,-8,4,7,18,42,47,30,17,35,34,56,40,52,53,67,59,57,85,52,64,65,62,57,55,46,51,79,53,63,76,42,65,64,39,55,57,56,54,50,43,44,36,38,49,26,24,26,5,-5,1,4,7,-0,-22,-7,-25,-6,-25,-35,-39,-49,-34,-38,-18,-50,-58,-71,-60,-62,-59,-65,-72,-81,-50,-66,-78,-53,-68,-83,-67,-64,-52,-52,-65,-63,-54,-56,-46,-56,-38,-37,-10,-34,-24,-7,-23,7,1,5,-7,1,10,-9,39,26,19,39,33,52,20,53,49,34,56,40,71,72,55,60,59,85,75,64,69,73,73,72,72,66,88,69,76,72,43,34,47,66,63,53,44,24,35,20,17,2,6,27,15,5,10,-1,-6,-8,-5,-20,-33,-12,-38,-28,-28,-41,-40,-55,-50,-56,-62,-43,-81,-59,-67,-47,-42,-72,-63,-61,-59,-64,-41,-46,-63,-55,-58,-71,-55,-49,-35,-59,-17,-72,-36,-5,-55,-32,-32,-24,-5,-16,7,-10,13,23,10,2,11,38,25,26,23,49,49,57,49,48,38,62,63,47,52,60,69,73,57,53,73,72,64,81,67,61,47,51,68,75,63,67,49,70,48,23,59,28,36,49,45,41,13,26,12,13,25,-5,-6,-35,-14,-10,-19,-39,-20,-25,-45,-46,-51,-57,-40,-48,-72,-58,-67,-39,-56,-47,-57,-66,-58,-62,-64,-88,-59,-84,-62,-41,-62,-51,-67,-29,-49,-35,-42,-59,-46,-32,-31,-45,-15,-28,10,6,-12,-2,8,4,6,24,27,18,32,31,39,34,56,63,38,25,47,46,55,75,75,75,61,69,76,79,43,67,63,56,82,50,68,48,47,78,61,46,57,26,66,30,26,14,39,28,12,22,27,20,28,1,20,-15,12,-20,27,-18,-34,-9,-20,-20,-17,-26,-40,-44,-54,-56,-64,-75,-59,-69,-66,-63,-66,-56,-78,-72,-56,-47,-78,-62,-69,-69,-51,-68,-53,-61,-63,-34,-40,-20,-40,-30,-36,-27,-7,-3,9,27,-31,13,11
--);

-- in=2000, out=2000, seno + ruído em freq 0,6(converge) (1)
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	-17,36,-19,26,18,9,65,12,53,36,22,65,25,70,44,35,82,25,64,52,46,92,30,79,59,46,85,29,77,49,34,92,27,76,51,28,84,17,59,38,11,59,-5,45,23,-3,48,-19,25,-3,-15,22,-41,-0,-26,-38,18,-54,-10,-41,-63,-11,-75,-20,-53,-73,-23,-88,-35,-60,-57,-34,-88,-42,-70,-78,-34,-87,-37,-59,-64,-25,-81,-32,-54,-54,-18,-69,-22,-29,-39,-3,-53,1,-22,-29,24,-37,27,-13,-1,27,-19,36,17,15,61,0,55,31,21,67,14,75,43,40,78,32,78,49,48,84,36,95,55,54,91,29,83,44,51,89,19,68,45,29,71,9,61,34,24,47,-3,53,10,-5,43,-23,27,1,-11,11,-42,6,-30,-32,-6,-52,-9,-35,-39,-17,-78,-25,-57,-63,-29,-83,-36,-65,-55,-28,-91,-37,-67,-61,-27,-95,-25,-56,-67,-28,-86,-28,-53,-53,-19,-74,-20,-44,-37,5,-58,8,-28,-14,11,-42,26,-19,-7,39,-16,45,19,14,52,-4,65,21,40,64,9,66,38,36,70,26,87,49,49,82,19,81,54,57,84,20,85,50,54,77,22,80,45,36,72,14,59,16,32,44,-6,57,10,5,39,-24,35,-13,2,9,-48,15,-24,-25,-2,-50,-7,-54,-39,-13,-76,-1,-63,-60,-31,-87,-37,-70,-70,-36,-71,-33,-84,-62,-39,-89,-32,-78,-61,-44,-95,-21,-60,-40,-27,-62,-2,-47,-35,-6,-61,-0,-45,-14,6,-36,30,-18,0,29,-14,47,3,15,41,-10,64,21,45,59,20,75,27,45,75,31,82,37,59,80,40,98,44,61,82,33,81,37,60,70,20,78,33,55,62,9,75,14,28,51,-7,53,11,20,29,-14,24,-17,-0,15,-33,19,-40,-16,-6,-59,3,-59,-31,-21,-74,-15,-71,-53,-27,-82,-20,-69,-58,-44,-82,-23,-83,-58,-52,-94,-33,-81,-52,-37,-74,-13,-62,-48,-22,-63,-17,-56,-17,-19,-54,6,-40,-7,8,-33,23,-17,0,24,-17,40,2,27,43,-10,71,16,27,57,11,75,29,63,76,29,83,39,59,69,28,87,42,62,76,36,81,40,58,68,25,81,27,52,54,25,78,16,39,37,-2,49,-0,16,28,-12,34,-20,-2,2,-32,12,-37,-13,-8,-53,4,-64,-28,-20,-71,-10,-71,-35,-46,-82,-29,-68,-53,-52,-78,-32,-88,-50,-40,-100,-21,-73,-25,-41,-81,-24,-71,-34,-38,-72,-12,-57,-24,-13,-50,4,-42,-11,-7,-22,26,-21,12,9,-21,48,-7,22,36,12,66,12,57,51,25,83,20,65,64,29,92,29,68,71,39,98,28,62,70,32,91,38,62,59,32,68,29,59,61,20,65,7,51,31,9,54,-4,34,28,-15,31,-17,11,4,-36,16,-49,-8,-20,-43,-2,-54,-27,-42,-67,-17,-81,-44,-38,-71,-24,-77,-53,-51,-84,-29,-85,-44,-51,-85,-29,-88,-36,-54,-77,-20,-83,-23,-41,-64,-10,-63,-9,-27,-53,14,-47,-5,-16,-29,33,-30,19,3,-20,44,-5,28,29,15,69,4,65,38,23,75,29,62,50,32,85,41,75,61,42,92,34,78,52,48,78,31,74,56,39,91,21,72,49,30,68,3,52,31,8,50,-3,37,19,3,31,-30,21,-2,-24,21,-47,6,-26,-48,5,-68,-11,-39,-54,-16,-65,-38,-50,-71,-26,-85,-37,-56,-77,-29,-83,-39,-57,-75,-18,-87,-39,-62,-72,-22,-79,-23,-42,-52,-19,-57,-15,-25,-37,10,-43,1,-17,-25,30,-31,17,4,-4,40,-13,47,24,13,60,6,59,39,22,91,13,80,43,38,86,12,69,52,49,86,33,80,54,44,90,30,78,58,43,81,19,70,42,31,64,5,50,25,2,55,0,29,12,-10,39,-39,16,-3,-19,19,-46,3,-34,-31,-3,-63,1,-50,-57,-16,-68,-25,-50,-67,-25,-77,-42,-68,-74,-40,-94,-43,-68,-64,-25,-87,-38,-64,-58,-28,-72,-15,-57,-54,-12,-67,-10,-23,-49,8,-51,6,-21,-3,15,-28,30,-11,-6,42,-13,42,7,24,47,6,64,41,37,75,24,85,50,42,78,28,99,44,46,79,26,85,55,53,80,26,77,42,47,78,26,80,28,29,62,5,56,20,16,51,-13,40,-2,7,30,-32,28,-15,-23,20,-49,6,-26,-30,-7,-59,-16,-48,-49,-25,-77,-24,-50,-74,-36,-75,-26,-70,-65,-33,-91,-32,-79,-59,-37,-84,-32,-53,-65,-20,-65,-23,-48,-54,-17,-59,-11,-47,-33,-3,-56,9,-28,-17,22,-40,36,-1,10,26,-4,46,10,26,59,9,67,29,40,60,21,87,31,51,73,30,89,41,56,80,26,81,35,56,82,37,82,42,55,75,25,81,36,43,58,6,67,21,22,39,-9,49,-6,12,19,-13,29,-29,-12,4,-50,0,-45,-25,-8,-55,-6,-58,-51,-19,-77,-29,-61,-55,-33,-86,-37,-64,-71,-43,-90,-30,-83,-55,-35,-86,-43,-73,-51,-32,-87,-13,-64,-37,-21,-62,2,-44,-23,-7,-38,5,-28,-8,10,-35,33,-5,15,29,-8,50,-0,25,39,9,72,15,38,68,22,74,32,63,84,31,80,42,61,84,34,86,42,61,87,24,83,32,56,71,24,80,36,54,57,3,64,7,22,45,-2,53,-9,5,11,-31,27,-19,-5,7,-45,10,-38,-26,-15,-56,-15,-61,-36,-22,-74,-15,-70,-56,-45,-77,-21,-79,-54,-47,-79,-33,-82,-60,-44,-79,-25,-79,-47,-43,-67,-20,-58,-33,-21,-55,-6,-54,-18,-18,-47,24,-40,-6,11,-28,38,-14,15,29,-2,50,6,34,43,16,65,24,55,63,31,75,35,61,59,48,89,36,74,74,30,76,38,70,71,32,87,38,60,67,19,76,25,52,55,13,68,6,34,31,-7,38,-18,12,11,-13,21,-38,-2,-2,-31,8,-54,-16,-20,-56,-1,-70,-28,-42,-66,-26,-79,-40,-53,-79,-25,-81,-40,-63,-84,-24,-99,-44,-45,-85,-27,-81,-41,-38,-76,-8,-77,-35,-31,-58,-4,-52,-17,-24,-50,17,-46,-6,6,-30,30,-12,20,30,-5,39,-5,47,43,7,60,17,49,54,25,83,21,70,64,43,93,29,76,74,40,83,38,78,61,46,90,34,64,63,16,83,24,62,45,21,61,-7,48,29,-4,46,-11,25,11,-14,33,-40,-6,-10,-35,13,-44,-8,-28,-61,-4,-71,-26,-39,-59,-13,-73,-31,-51,-74,-33,-75,-46,-55,-71,-30,-82,-42,-55,-75,-31,-91,-39,-41,-63,-14,-77,-21,-28,-66,-8,-57,-7,-13,-46,19,-36,13,-1,-10,34,-35,27,20,-5,53,-5,42,29,13,65,13,63,53,33,82,21,74,59,33,89,26,85,63,50,90,41,81,62,38,83,37,73,53,33,67,15,58,37,25,68,5,47,25,15,46,-13,27,7,-24,30,-27,17,-24,-35,14,-51,-2,-36,-45,-9,-65,-16,-46,-60,-16,-86,-33,-50,-65,-34,-89,-36,-56,-77,-37,-88,-39,-64,-74,-28,-90,-49,-54,-56,-8,-84,-23,-48,-41,-9,-62,-2,-19,-33,16,-45,5,-14,-13,25,-21,38,9,8,53,-10,51,30,21,62,20,66,41,46,71,17,68,43,50,73,33,87,56,38,91,38,87,51,47,86,40,80,53,34,76,12,70,25,23,56,1,65,15,19,42,-7,25,-5,-5,30,-30,16,-24,-25,8,-58,3,-39,-31,-3,-64,-21,-64,-55,-27,-74,-21,-74,-68,-29,-90,-44,-58,-66,-31,-93,-27,-60,-67,-38,-86,-26,-64,-64,-11,-74,-15,-58,-45,-6,-67,3,-26,-28,10,-45,16,-17,-4,30,-23,32,13,17,47,-2,50,23,26,63,16,72,36,39,73,24,79,45,50,84,21,98,53,49,87,20,81,49,56,81,34,83,37,38,68,13,74,35,29,61,8,65,21,8,43,-8,30,-4,5,23,-39,18,-25,-17,7,-58,10,-50,-35,-11,-60,-17,-52,-59,-29,-74,-20,-64,-59,-33,-90,-29,-82,-65,-38,-86,-49,-71,-65,-40,-74,-27,-60,-51,-24,-75,-19,-63,-38,-15,-71,-2,-50,-23,7,-46,20,-13,-2,14,-27,34,-4,23,49,-6,47,13,28,62,7,72,29,51,70,22,93,34,55,77,28,84,38,50,72,37,83,41,63,67,29,86,27,50,69,20,76,26,40,57,5,62,18,24,39,-8,38,-15,4,20,-26,26,-33,-9,-2,-42,6,-48,-32,-22,-63,-8,-48,-44,-34,-86,-24,-74,-53,-42,-91,-37,-72,-59,-50,-83,-32,-88,-58,-43,-81,-22,-77,-53,-35,-78,-14,-68,-35,-20,-50,-2,-45,-13,-6,-34,23,-23,-4,14,-23,28,1,22,31,0,56,16,28,55,13,65,26,45,70,30,80,33,59,81,36,89,40,68,77,36,93,38,75,74,36,91,25,47,60,28,82,24,46,43,7,55,-0,19,26,-6,44,-15,14,13,-30,24,-29,-9,-11,-42,1,-49,-21,-24,-62,-15,-67,-41,-41,-70,-33,-77,-51,-39,-74,-32,-82,-51,-46,-85,-19,-75,-51,-44,-81,-31,-77,-41,-31,-77,-1,-79,-29,-11,-68,-1,-53,-15,-3,-41,26,-34,11,19,-20,33,-15,32,28,-3,52,11,47,52,16,72,13,60,61,22,80,29,69,70,31,84,38,73,68,43,91,32,62,60,36,93,30,68,55,33,75,7,58,39,10,69,9,42,24,-2,43,-15,26,6,-26,12,-37,1,-10,-50,9,-51,-23,-31,-64,-16,-66,-32,-51,-74,-27,-71,-41,-44,-77,-30,-83,-46,-54,-93,-27,-96,-45,-43,-79,-21,-85,-26,-43,-62,-13,-76,-28,-30,-54,-7,-49,-12,-2,-28,17,-34,14,4,-18,43,-11,28,26,3,59,1,55,49,15,60,14,58,52,38,89,33,70,63,43,95,21,76,61,36,97,25,77,53,30,93,27,64,53,17,83,7,49,27,16,58,-9,39,25,-1,50,-23,30,-4,-13,18,-20,3,-22,-32,8,-51,-5,-28,-55,-10,-74,-30,-53,-77,-24,-87,-40,-57,-77,-26,-94,-45,-56,-69,-37,-88,-43,-62,-70,-31,-81,-36,-55,-57,-13,-61,-20,-34,-51,-0,-47,5,-9,-14,6,-29,1
--);

-- in=2000, out=2000, seno freq 0,01 + ruído em freq 0,6(converge) (1)
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	-17,36,-19,26,18,9,65,12,53,36,22,65,25,70,44,35,82,25,64,52,46,92,30,79,59,46,85,29,77,49,34,92,27,76,51,28,84,17,59,38,11,59,-5,45,23,-3,48,-19,25,-3,-15,22,-41,-0,-26,-38,18,-54,-10,-41,-63,-11,-75,-20,-53,-73,-23,-88,-35,-60,-57,-34,-88,-42,-70,-78,-34,-87,-37,-59,-64,-25,-81,-32,-54,-54,-18,-69,-22,-29,-39,-3,-53,1,-22,-29,24,-37,27,-13,-1,27,-19,36,17,15,61,0,55,31,21,67,14,75,43,40,78,32,78,49,48,84,36,95,55,54,91,29,83,44,51,89,19,68,45,29,71,9,61,34,24,47,-3,53,10,-5,43,-23,27,1,-11,11,-42,6,-30,-32,-6,-52,-9,-35,-39,-17,-78,-25,-57,-63,-29,-83,-36,-65,-55,-28,-91,-37,-67,-61,-27,-95,-25,-56,-67,-28,-86,-28,-53,-53,-19,-74,-20,-44,-37,5,-58,8,-28,-14,11,-42,26,-19,-7,39,-16,45,19,14,52,-4,65,21,40,64,9,66,38,36,70,26,87,49,49,82,19,81,54,57,84,20,85,50,54,77,22,80,45,36,72,14,59,16,32,44,-6,57,10,5,39,-24,35,-13,2,9,-48,15,-24,-25,-2,-50,-7,-54,-39,-13,-76,-1,-63,-60,-31,-87,-37,-70,-70,-36,-71,-33,-84,-62,-39,-89,-32,-78,-61,-44,-95,-21,-60,-40,-27,-62,-2,-47,-35,-6,-61,-0,-45,-14,6,-36,30,-18,0,29,-14,47,3,15,41,-10,64,21,45,59,20,75,27,45,75,31,82,37,59,80,40,98,44,61,82,33,81,37,60,70,20,78,33,55,62,9,75,14,28,51,-7,53,11,20,29,-14,24,-17,-0,15,-33,19,-40,-16,-6,-59,3,-59,-31,-21,-74,-15,-71,-53,-27,-82,-20,-69,-58,-44,-82,-23,-83,-58,-52,-94,-33,-81,-52,-37,-74,-13,-62,-48,-22,-63,-17,-56,-17,-19,-54,6,-40,-7,8,-33,23,-17,0,24,-17,40,2,27,43,-10,71,16,27,57,11,75,29,63,76,29,83,39,59,69,28,87,42,62,76,36,81,40,58,68,25,81,27,52,54,25,78,16,39,37,-2,49,-0,16,28,-12,34,-20,-2,2,-32,12,-37,-13,-8,-53,4,-64,-28,-20,-71,-10,-71,-35,-46,-82,-29,-68,-53,-52,-78,-32,-88,-50,-40,-100,-21,-73,-25,-41,-81,-24,-71,-34,-38,-72,-12,-57,-24,-13,-50,4,-42,-11,-7,-22,26,-21,12,9,-21,48,-7,22,36,12,66,12,57,51,25,83,20,65,64,29,92,29,68,71,39,98,28,62,70,32,91,38,62,59,32,68,29,59,61,20,65,7,51,31,9,54,-4,34,28,-15,31,-17,11,4,-36,16,-49,-8,-20,-43,-2,-54,-27,-42,-67,-17,-81,-44,-38,-71,-24,-77,-53,-51,-84,-29,-85,-44,-51,-85,-29,-88,-36,-54,-77,-20,-83,-23,-41,-64,-10,-63,-9,-27,-53,14,-47,-5,-16,-29,33,-30,19,3,-20,44,-5,28,29,15,69,4,65,38,23,75,29,62,50,32,85,41,75,61,42,92,34,78,52,48,78,31,74,56,39,91,21,72,49,30,68,3,52,31,8,50,-3,37,19,3,31,-30,21,-2,-24,21,-47,6,-26,-48,5,-68,-11,-39,-54,-16,-65,-38,-50,-71,-26,-85,-37,-56,-77,-29,-83,-39,-57,-75,-18,-87,-39,-62,-72,-22,-79,-23,-42,-52,-19,-57,-15,-25,-37,10,-43,1,-17,-25,30,-31,17,4,-4,40,-13,47,24,13,60,6,59,39,22,91,13,80,43,38,86,12,69,52,49,86,33,80,54,44,90,30,78,58,43,81,19,70,42,31,64,5,50,25,2,55,0,29,12,-10,39,-39,16,-3,-19,19,-46,3,-34,-31,-3,-63,1,-50,-57,-16,-68,-25,-50,-67,-25,-77,-42,-68,-74,-40,-94,-43,-68,-64,-25,-87,-38,-64,-58,-28,-72,-15,-57,-54,-12,-67,-10,-23,-49,8,-51,6,-21,-3,15,-28,30,-11,-6,42,-13,42,7,24,47,6,64,41,37,75,24,85,50,42,78,28,99,44,46,79,26,85,55,53,80,26,77,42,47,78,26,80,28,29,62,5,56,20,16,51,-13,40,-2,7,30,-32,28,-15,-23,20,-49,6,-26,-30,-7,-59,-16,-48,-49,-25,-77,-24,-50,-74,-36,-75,-26,-70,-65,-33,-91,-32,-79,-59,-37,-84,-32,-53,-65,-20,-65,-23,-48,-54,-17,-59,-11,-47,-33,-3,-56,9,-28,-17,22,-40,36,-1,10,26,-4,46,10,26,59,9,67,29,40,60,21,87,31,51,73,30,89,41,56,80,26,81,35,56,82,37,82,42,55,75,25,81,36,43,58,6,67,21,22,39,-9,49,-6,12,19,-13,29,-29,-12,4,-50,0,-45,-25,-8,-55,-6,-58,-51,-19,-77,-29,-61,-55,-33,-86,-37,-64,-71,-43,-90,-30,-83,-55,-35,-86,-43,-73,-51,-32,-87,-13,-64,-37,-21,-62,2,-44,-23,-7,-38,5,-28,-8,10,-35,33,-5,15,29,-8,50,-0,25,39,9,72,15,38,68,22,74,32,63,84,31,80,42,61,84,34,86,42,61,87,24,83,32,56,71,24,80,36,54,57,3,64,7,22,45,-2,53,-9,5,11,-31,27,-19,-5,7,-45,10,-38,-26,-15,-56,-15,-61,-36,-22,-74,-15,-70,-56,-45,-77,-21,-79,-54,-47,-79,-33,-82,-60,-44,-79,-25,-79,-47,-43,-67,-20,-58,-33,-21,-55,-6,-54,-18,-18,-47,24,-40,-6,11,-28,38,-14,15,29,-2,50,6,34,43,16,65,24,55,63,31,75,35,61,59,48,89,36,74,74,30,76,38,70,71,32,87,38,60,67,19,76,25,52,55,13,68,6,34,31,-7,38,-18,12,11,-13,21,-38,-2,-2,-31,8,-54,-16,-20,-56,-1,-70,-28,-42,-66,-26,-79,-40,-53,-79,-25,-81,-40,-63,-84,-24,-99,-44,-45,-85,-27,-81,-41,-38,-76,-8,-77,-35,-31,-58,-4,-52,-17,-24,-50,17,-46,-6,6,-30,30,-12,20,30,-5,39,-5,47,43,7,60,17,49,54,25,83,21,70,64,43,93,29,76,74,40,83,38,78,61,46,90,34,64,63,16,83,24,62,45,21,61,-7,48,29,-4,46,-11,25,11,-14,33,-40,-6,-10,-35,13,-44,-8,-28,-61,-4,-71,-26,-39,-59,-13,-73,-31,-51,-74,-33,-75,-46,-55,-71,-30,-82,-42,-55,-75,-31,-91,-39,-41,-63,-14,-77,-21,-28,-66,-8,-57,-7,-13,-46,19,-36,13,-1,-10,34,-35,27,20,-5,53,-5,42,29,13,65,13,63,53,33,82,21,74,59,33,89,26,85,63,50,90,41,81,62,38,83,37,73,53,33,67,15,58,37,25,68,5,47,25,15,46,-13,27,7,-24,30,-27,17,-24,-35,14,-51,-2,-36,-45,-9,-65,-16,-46,-60,-16,-86,-33,-50,-65,-34,-89,-36,-56,-77,-37,-88,-39,-64,-74,-28,-90,-49,-54,-56,-8,-84,-23,-48,-41,-9,-62,-2,-19,-33,16,-45,5,-14,-13,25,-21,38,9,8,53,-10,51,30,21,62,20,66,41,46,71,17,68,43,50,73,33,87,56,38,91,38,87,51,47,86,40,80,53,34,76,12,70,25,23,56,1,65,15,19,42,-7,25,-5,-5,30,-30,16,-24,-25,8,-58,3,-39,-31,-3,-64,-21,-64,-55,-27,-74,-21,-74,-68,-29,-90,-44,-58,-66,-31,-93,-27,-60,-67,-38,-86,-26,-64,-64,-11,-74,-15,-58,-45,-6,-67,3,-26,-28,10,-45,16,-17,-4,30,-23,32,13,17,47,-2,50,23,26,63,16,72,36,39,73,24,79,45,50,84,21,98,53,49,87,20,81,49,56,81,34,83,37,38,68,13,74,35,29,61,8,65,21,8,43,-8,30,-4,5,23,-39,18,-25,-17,7,-58,10,-50,-35,-11,-60,-17,-52,-59,-29,-74,-20,-64,-59,-33,-90,-29,-82,-65,-38,-86,-49,-71,-65,-40,-74,-27,-60,-51,-24,-75,-19,-63,-38,-15,-71,-2,-50,-23,7,-46,20,-13,-2,14,-27,34,-4,23,49,-6,47,13,28,62,7,72,29,51,70,22,93,34,55,77,28,84,38,50,72,37,83,41,63,67,29,86,27,50,69,20,76,26,40,57,5,62,18,24,39,-8,38,-15,4,20,-26,26,-33,-9,-2,-42,6,-48,-32,-22,-63,-8,-48,-44,-34,-86,-24,-74,-53,-42,-91,-37,-72,-59,-50,-83,-32,-88,-58,-43,-81,-22,-77,-53,-35,-78,-14,-68,-35,-20,-50,-2,-45,-13,-6,-34,23,-23,-4,14,-23,28,1,22,31,0,56,16,28,55,13,65,26,45,70,30,80,33,59,81,36,89,40,68,77,36,93,38,75,74,36,91,25,47,60,28,82,24,46,43,7,55,-0,19,26,-6,44,-15,14,13,-30,24,-29,-9,-11,-42,1,-49,-21,-24,-62,-15,-67,-41,-41,-70,-33,-77,-51,-39,-74,-32,-82,-51,-46,-85,-19,-75,-51,-44,-81,-31,-77,-41,-31,-77,-1,-79,-29,-11,-68,-1,-53,-15,-3,-41,26,-34,11,19,-20,33,-15,32,28,-3,52,11,47,52,16,72,13,60,61,22,80,29,69,70,31,84,38,73,68,43,91,32,62,60,36,93,30,68,55,33,75,7,58,39,10,69,9,42,24,-2,43,-15,26,6,-26,12,-37,1,-10,-50,9,-51,-23,-31,-64,-16,-66,-32,-51,-74,-27,-71,-41,-44,-77,-30,-83,-46,-54,-93,-27,-96,-45,-43,-79,-21,-85,-26,-43,-62,-13,-76,-28,-30,-54,-7,-49,-12,-2,-28,17,-34,14,4,-18,43,-11,28,26,3,59,1,55,49,15,60,14,58,52,38,89,33,70,63,43,95,21,76,61,36,97,25,77,53,30,93,27,64,53,17,83,7,49,27,16,58,-9,39,25,-1,50,-23,30,-4,-13,18,-20,3,-22,-32,8,-51,-5,-28,-55,-10,-74,-30,-53,-77,-24,-87,-40,-57,-77,-26,-94,-45,-56,-69,-37,-88,-43,-62,-70,-31,-81,-36,-55,-57,-13,-61,-20,-34,-51,-0,-47,5,-9,-14,6,-29,1
--);
	
-- in=2000, out=2000, seno freq 0,01  + ruído aleatório (white gaussian noise) (converge mais ou menos)
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	-2,9,9,2,20,34,51,57,40,43,45,36,71,62,46,59,59,59,38,55,75,75,65,67,66,71,59,64,63,48,50,80,67,67,62,45,74,57,43,50,24,35,26,30,36,11,32,15,6,-1,5,-4,-12,-28,-28,-26,8,-22,-30,-42,-63,-40,-51,-38,-55,-71,-52,-66,-60,-60,-30,-68,-62,-71,-76,-73,-68,-58,-63,-56,-49,-54,-54,-60,-53,-36,-48,-40,-54,-12,-20,-34,-22,-20,-16,-19,8,-7,14,-15,22,-5,13,14,30,37,48,35,36,44,32,45,49,64,56,58,57,76,59,59,67,63,80,91,71,78,76,66,66,51,75,79,51,41,61,36,52,40,40,53,41,17,32,39,20,-4,27,8,2,20,1,-22,-14,-23,-26,-25,-40,-16,-39,-18,-23,-46,-56,-57,-51,-61,-59,-54,-70,-57,-36,-50,-66,-69,-57,-49,-46,-76,-45,-38,-66,-54,-63,-60,-39,-46,-45,-50,-55,-32,-27,-8,-32,-13,-16,3,-12,-17,6,-15,-2,27,21,28,48,23,36,28,51,35,61,47,39,37,57,39,46,63,72,73,58,66,42,53,79,73,69,45,63,75,70,59,56,61,73,40,61,51,28,26,45,17,25,42,31,5,25,4,12,2,17,-19,-28,-12,-2,-21,-23,-13,-41,-48,-34,-29,-53,-13,-51,-68,-55,-64,-81,-58,-82,-58,-25,-66,-84,-62,-64,-64,-66,-73,-65,-80,-83,-50,-43,-31,-52,-24,-22,-27,-34,-23,-39,-37,-40,-8,-15,-4,10,-1,1,15,24,27,25,13,23,13,44,46,60,44,60,52,45,45,68,73,56,56,67,71,85,85,70,68,74,71,50,58,69,54,50,50,57,67,49,37,57,31,24,41,19,26,44,23,12,21,-16,2,-0,3,2,-8,-26,-14,-22,-37,-24,-48,-30,-37,-52,-47,-59,-65,-36,-58,-46,-45,-68,-65,-52,-48,-72,-67,-82,-78,-72,-70,-58,-53,-43,-36,-37,-59,-31,-30,-58,-37,-8,-40,-28,-25,-20,-6,-0,-2,-8,10,-11,15,12,7,33,27,36,7,57,44,8,51,36,48,59,73,80,64,55,72,54,57,56,59,74,57,72,73,48,72,52,61,54,55,55,48,42,65,62,45,34,22,24,15,28,2,22,20,3,5,-17,-13,-3,-26,-11,-22,-15,-29,-23,-51,-37,-24,-52,-38,-50,-40,-67,-65,-68,-35,-70,-71,-51,-70,-73,-60,-44,-98,-47,-44,-12,-51,-63,-62,-47,-42,-54,-56,-47,-31,-35,-16,-25,-32,-15,-26,-20,16,-4,11,3,-5,-2,25,21,5,35,50,46,44,62,50,61,66,48,66,67,57,76,58,63,75,72,82,51,45,70,56,69,75,50,53,61,26,67,52,69,48,33,32,48,20,40,25,26,30,34,5,-3,19,-2,2,-20,-17,-31,-23,-30,-15,-37,-23,-46,-59,-52,-53,-65,-71,-38,-49,-57,-48,-82,-57,-70,-63,-60,-61,-56,-74,-63,-68,-47,-66,-63,-51,-66,-30,-49,-47,-43,-37,-13,-33,-40,-7,-20,-24,-27,-7,14,-1,8,-6,-9,18,32,6,32,47,53,34,69,35,48,51,72,48,48,55,61,90,67,66,70,71,71,68,46,82,42,68,64,59,67,77,54,69,55,59,42,29,38,33,28,20,33,25,26,36,-1,-6,10,1,-4,-4,-21,-3,-30,-36,-19,-48,-24,-41,-33,-48,-26,-68,-51,-58,-58,-60,-58,-56,-66,-60,-51,-60,-55,-61,-36,-62,-64,-70,-61,-52,-54,-39,-37,-29,-58,-19,-36,-16,-14,-13,-6,-20,-16,-7,12,-1,-6,9,17,14,18,37,35,34,39,42,46,50,37,89,43,77,47,57,69,31,43,58,75,62,71,63,61,63,74,68,62,76,66,60,52,54,51,51,37,36,25,32,5,34,43,-3,23,-3,19,-22,-12,10,-3,-3,-18,-21,-37,-11,-32,-34,-7,-53,-52,-43,-32,-50,-40,-62,-51,-40,-77,-69,-70,-78,-72,-77,-67,-47,-46,-59,-71,-63,-41,-59,-36,-30,-57,-45,-36,-39,-35,1,-51,-11,-22,-18,-12,29,-15,9,14,-9,1,24,20,19,9,45,17,44,48,67,58,60,67,80,74,54,57,67,100,54,57,55,57,66,76,71,57,60,51,53,63,60,68,68,34,35,40,35,30,32,22,32,15,13,4,21,6,-6,6,-4,-23,5,-22,-22,-7,-21,-33,-27,-51,-38,-45,-57,-52,-55,-26,-87,-67,-36,-50,-61,-62,-55,-67,-60,-80,-49,-65,-54,-64,-27,-70,-35,-20,-54,-27,-57,-41,-21,-43,-38,-29,-26,-31,-19,-14,-14,9,-18,20,23,25,-2,40,21,28,38,50,51,48,53,52,38,60,78,45,62,54,70,71,58,65,65,57,52,44,65,71,81,56,65,67,63,64,64,62,53,38,36,46,45,23,16,21,26,7,20,-10,33,3,-24,-12,-21,-29,-40,-38,-22,-27,-20,-36,-48,-62,-34,-53,-72,-40,-60,-54,-63,-80,-37,-88,-68,-67,-61,-76,-53,-50,-59,-94,-59,-50,-51,-72,-38,-49,-32,-39,-30,-19,-20,-18,-25,4,-32,-4,-7,-7,-8,9,25,23,15,30,26,17,25,17,46,54,32,36,64,59,44,58,76,88,68,49,72,64,83,70,58,69,63,92,49,55,52,56,64,58,56,72,64,46,25,37,24,10,37,32,30,10,-10,-15,-12,-6,8,-12,-3,-21,-23,-12,-38,-32,-28,-59,-45,-42,-31,-51,-46,-49,-73,-68,-48,-48,-61,-64,-66,-48,-71,-64,-77,-59,-49,-58,-63,-54,-63,-32,-56,-26,-36,-29,-21,-39,-33,-20,-38,-21,8,-20,-13,6,1,19,16,12,25,38,23,39,31,37,58,38,62,59,65,75,45,72,60,47,99,67,67,81,72,57,34,69,71,68,62,61,75,53,67,40,46,56,47,52,41,43,31,24,18,15,-5,-2,-7,-6,21,-21,-25,-17,-13,2,-29,-40,-28,-31,-34,-30,-56,-38,-63,-40,-69,-61,-52,-74,-60,-58,-58,-46,-88,-66,-53,-94,-53,-49,-69,-61,-58,-54,-41,-58,-30,-59,-51,-36,-33,-34,-20,-29,-39,-32,-7,-25,-26,9,-10,2,29,11,42,24,1,25,49,50,31,27,53,35,58,54,64,50,67,68,81,75,59,73,84,71,51,77,75,58,85,67,71,49,69,25,63,61,56,43,49,29,9,41,26,12,15,19,10,7,9,6,-24,-37,-18,-16,-17,-13,-24,-38,-54,-36,-53,-45,-44,-35,-39,-44,-45,-57,-57,-74,-40,-70,-59,-46,-64,-51,-61,-58,-56,-69,-75,-59,-35,-39,-40,-53,-33,-19,-60,-42,-26,-19,-1,-34,-1,1,6,6,24,12,-15,16,33,14,34,28,27,33,33,42,51,56,68,62,63,54,65,71,49,70,58,82,74,82,68,86,72,72,58,55,82,60,60,52,31,45,36,38,49,46,39,29,29,43,18,18,2,9,-21,4,8,2,-36,-27,-11,-23,-19,-41,-29,-43,-35,-33,-47,-46,-43,-68,-58,-43,-49,-71,-65,-59,-49,-68,-75,-60,-64,-67,-65,-58,-69,-90,-50,-34,-24,-65,-47,-48,-16,-38,-34,-17,-3,-14,-1,-15,-21,-9,8,-2,19,30,21,33,38,22,39,48,40,41,69,52,56,79,46,50,44,50,76,40,76,76,70,44,77,83,75,62,65,68,93,66,72,43,55,40,54,24,32,26,32,59,21,40,14,32,-9,-3,7,8,3,-10,-25,-16,-19,-37,-19,-36,-11,-23,-32,-53,-75,-47,-60,-41,-41,-82,-65,-55,-66,-84,-42,-56,-56,-71,-46,-45,-61,-73,-60,-50,-59,-62,-22,-42,-36,-57,-34,-24,-42,-14,-5,-15,-8,-13,-5,-3,16,17,14,10,42,41,33,40,27,45,40,50,62,58,57,53,57,65,59,64,65,72,48,94,76,57,75,44,55,69,72,65,78,63,49,41,45,42,56,57,33,44,46,52,44,3,23,31,-7,9,16,1,-18,-14,-14,-12,-13,-40,-10,-49,-33,-34,-25,-52,-36,-69,-58,-41,-46,-49,-59,-55,-67,-58,-82,-68,-62,-56,-100,-57,-69,-68,-34,-58,-39,-47,-42,-46,-51,-57,-32,-36,-53,-30,-44,-16,-6,-17,-1,17,9,-8,4,7,18,42,47,30,17,35,34,56,40,52,53,67,59,57,85,52,64,65,62,57,55,46,51,79,53,63,76,42,65,64,39,55,57,56,54,50,43,44,36,38,49,26,24,26,5,-5,1,4,7,-0,-22,-7,-25,-6,-25,-35,-39,-49,-34,-38,-18,-50,-58,-71,-60,-62,-59,-65,-72,-81,-50,-66,-78,-53,-68,-83,-67,-64,-52,-52,-65,-63,-54,-56,-46,-56,-38,-37,-10,-34,-24,-7,-23,7,1,5,-7,1,10,-9,39,26,19,39,33,52,20,53,49,34,56,40,71,72,55,60,59,85,75,64,69,73,73,72,72,66,88,69,76,72,43,34,47,66,63,53,44,24,35,20,17,2,6,27,15,5,10,-1,-6,-8,-5,-20,-33,-12,-38,-28,-28,-41,-40,-55,-50,-56,-62,-43,-81,-59,-67,-47,-42,-72,-63,-61,-59,-64,-41,-46,-63,-55,-58,-71,-55,-49,-35,-59,-17,-72,-36,-5,-55,-32,-32,-24,-5,-16,7,-10,13,23,10,2,11,38,25,26,23,49,49,57,49,48,38,62,63,47,52,60,69,73,57,53,73,72,64,81,67,61,47,51,68,75,63,67,49,70,48,23,59,28,36,49,45,41,13,26,12,13,25,-5,-6,-35,-14,-10,-19,-39,-20,-25,-45,-46,-51,-57,-40,-48,-72,-58,-67,-39,-56,-47,-57,-66,-58,-62,-64,-88,-59,-84,-62,-41,-62,-51,-67,-29,-49,-35,-42,-59,-46,-32,-31,-45,-15,-28,10,6,-12,-2,8,4,6,24,27,18,32,31,39,34,56,63,38,25,47,46,55,75,75,75,61,69,76,79,43,67,63,56,82,50,68,48,47,78,61,46,57,26,66,30,26,14,39,28,12,22,27,20,28,1,20,-15,12,-20,27,-18,-34,-9,-20,-20,-17,-26,-40,-44,-54,-56,-64,-75,-59,-69,-66,-63,-66,-56,-78,-72,-56,-47,-78,-62,-69,-69,-51,-68,-53,-61,-63,-34,-40,-20,-40,-30,-36,-27,-7,-3,9,27,-31,13,11
--);

 --in=2000, out=2000, seno freq 0,01  + ruído em freq 0.6,0.7 e 0.8 (não converge)
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	-264,102,127,96,90,8,19,4,349,83,-114,246,217,211,180,130,161,69,471,204,-93,289,220,305,182,131,202,104,464,215,-42,283,251,204,164,138,108,49,377,124,-135,244,118,149,31,-46,28,-81,248,14,-291,44,-25,58,-87,-145,-84,-184,202,-83,-399,-31,-153,-51,-157,-224,-226,-237,105,-196,-445,-156,-191,-149,-253,-288,-212,-307,78,-234,-466,-72,-142,-104,-165,-187,-191,-174,107,-155,-333,-28,-70,-71,-88,-64,-20,-149,210,15,-231,118,27,132,59,17,38,50,371,91,-143,244,170,189,176,130,123,126,449,181,-40,275,276,279,234,95,156,155,483,191,-41,287,214,227,158,68,107,19,435,116,-198,169,96,126,44,-8,41,-116,260,14,-291,63,18,20,-55,-137,-97,-197,164,-129,-310,-39,-165,-70,-171,-233,-197,-321,37,-157,-409,-87,-162,-152,-204,-314,-229,-358,95,-224,-436,-71,-147,-76,-203,-204,-167,-275,105,-85,-393,12,-68,-20,-90,-90,-38,-127,202,15,-294,106,100,115,77,-29,90,3,335,110,-122,283,189,197,165,172,149,122,461,189,-10,315,236,281,226,166,215,80,476,216,-33,306,209,207,155,119,129,74,369,70,-187,179,101,155,67,-4,-23,-102,279,-39,-251,91,-4,47,-36,-111,-87,-232,112,-70,-389,-3,-140,-61,-194,-192,-203,-324,19,-204,-412,-50,-182,-115,-258,-252,-268,-309,71,-230,-472,-98,-159,-112,-165,-177,-173,-237,164,-141,-338,16,-72,33,-13,-111,-53,-144,210,-25,-190,105,78,137,48,21,60,-24,287,142,-126,268,186,234,136,125,179,49,387,237,-78,295,256,273,158,147,153,116,433,223,-18,284,204,239,181,64,114,12,364,176,-174,202,137,81,67,45,-8,-103,289,-82,-256,84,-2,-4,-30,-134,-84,-195,161,-120,-386,-38,-68,-84,-181,-221,-176,-270,93,-178,-432,-79,-190,-93,-197,-313,-234,-279,27,-188,-450,-144,-224,-135,-146,-243,-152,-264,116,-128,-324,-25,-79,-29,-50,-110,-51,-134,209,-33,-229,124,88,78,39,15,102,15,352,144,-124,222,195,182,165,111,177,17,472,174,-61,349,267,287,227,164,180,100,474,208,-62,312,247,237,173,96,102,74,390,111,-136,220,150,137,58,-70,26,-64,302,-42,-222,41,-7,29,-33,-135,-80,-170,128,-133,-444,23,-170,-75,-119,-240,-216,-246,83,-176,-428,-87,-242,-154,-225,-221,-230,-226,23,-227,-429,-81,-169,-79,-176,-212,-115,-265,145,-130,-385,56,-27,-36,-75,-53,-71,-101,250,19,-228,192,75,134,74,14,68,16,319,112,-99,190,185,228,194,116,183,64,449,208,-29,289,280,272,184,108,165,159,471,166,-105,262,223,212,178,103,126,32,397,135,-173,116,101,123,38,11,33,-28,293,-26,-226,72,20,8,-6,-164,-114,-213,139,-164,-376,-83,-166,-76,-165,-213,-212,-289,70,-207,-462,-105,-179,-119,-205,-246,-191,-284,33,-157,-480,-148,-134,-101,-153,-227,-151,-244,125,-162,-323,12,-11,-12,-85,-71,-71,-182,238,24,-234,128,54,140,45,-11,71,-31,379,84,-117,251,170,231,243,121,192,54,444,210,-91,291,238,301,213,116,170,88,503,158,-90,313,218,230,184,112,164,-18,382,148,-116,144,86,94,78,-14,-62,-89,284,44,-275,119,42,64,-72,-179,-131,-208,169,-153,-405,-72,-74,-105,-124,-179,-174,-291,45,-193,-447,-86,-209,-139,-231,-223,-183,-349,73,-157,-471,-48,-171,-115,-125,-169,-124,-222,114,-143,-354,-33,-78,-33,-72,-90,-67,-104,265,-45,-232,129,103,55,28,53,70,24,376,106,-155,265,134,175,197,166,151,132,498,240,-125,246,246,255,191,83,198,103,461,158,-99,286,196,287,160,88,140,36,399,127,-189,209,137,165,37,23,32,-37,290,5,-245,74,-49,0,-42,-159,-93,-200,172,-100,-365,-35,-139,-47,-176,-234,-202,-324,70,-212,-475,-120,-176,-103,-214,-295,-246,-215,41,-187,-438,-59,-78,-110,-202,-248,-151,-228,155,-75,-394,38,-23,-1,-63,-133,-96,-102,269,1,-247,180,50,130,98,85,7,26,375,126,-156,280,135,254,173,88,165,51,419,201,-28,339,257,246,222,128,179,94,399,220,-56,274,201,227,145,106,173,97,379,102,-190,204,91,122,57,-34,30,-98,249,26,-312,59,-32,40,-67,-162,-119,-233,143,-125,-348,-105,-90,-64,-166,-232,-239,-293,59,-122,-446,-79,-201,-154,-245,-312,-214,-285,11,-210,-500,-108,-157,-107,-131,-258,-147,-168,134,-135,-351,-6,-115,-53,-76,-126,-69,-162,229,-31,-252,97,35,134,102,-20,77,-8,348,159,-124,255,164,212,178,81,146,139,474,260,-87,302,197,289,178,164,164,93,464,156,-61,268,170,253,228,110,175,41,394,88,-135,184,144,138,100,-16,50,-94,276,16,-255,80,-16,59,-7,-100,-74,-196,134,-138,-379,-63,-149,-76,-191,-202,-200,-244,69,-197,-430,-102,-188,-134,-188,-212,-220,-328,69,-179,-443,-48,-104,-81,-194,-193,-246,-225,137,-107,-457,-61,-38,-48,-36,-115,-31,-109,202,20,-255,118,54,54,51,34,69,3,373,142,-99,239,143,238,243,176,150,32,447,170,-9,261,171,288,191,181,174,61,451,201,-80,322,181,265,152,84,201,70,397,96,-162,186,99,129,40,19,16,-112,268,-11,-281,95,-26,54,-59,-145,-70,-185,104,-169,-339,-32,-104,-115,-185,-258,-224,-279,71,-199,-427,-113,-227,-149,-159,-229,-252,-274,25,-226,-463,-50,-177,-111,-110,-143,-186,-226,108,-83,-373,-16,-71,37,-77,-93,-100,-85,289,27,-229,183,50,110,70,12,55,-22,372,148,-136,272,151,243,176,151,235,90,445,160,-68,293,210,320,195,189,192,144,462,199,-90,267,251,256,206,125,139,28,339,104,-157,172,135,132,55,-15,44,-86,281,36,-244,52,-85,6,-74,-136,-97,-203,168,-87,-407,-58,-105,-124,-143,-219,-206,-261,11,-216,-470,-155,-144,-151,-131,-261,-258,-287,49,-240,-453,-111,-99,-158,-96,-192,-170,-188,102,-130,-344,22,-20,-4,-126,-114,-52,-144,218,-6,-242,103,70,108,67,59,108,-13,402,137,-106,293,129,216,190,84,124,66,414,240,-58,333,182,222,246,211,158,129,448,170,-96,278,201,240,194,106,113,35,405,103,-167,232,100,146,21,29,-1,-48,272,-6,-259,24,-12,-13,-38,-117,-92,-194,149,-134,-385,-19,-76,-85,-138,-182,-228,-294,100,-170,-471,-131,-168,-146,-177,-286,-220,-258,88,-251,-417,-82,-158,-111,-167,-205,-201,-289,80,-183,-355,37,-94,38,-59,-88,-31,-123,248,-50,-292,113,82,105,64,-1,1,8,347,109,-106,266,205,160,176,177,155,80,401,230,-79,313,173,254,232,120,199,139,467,189,-70,250,231,250,191,102,99,36,337,127,-115,238,146,181,34,44,20,-57,240,18,-230,49,52,-16,-30,-144,-133,-164,132,-120,-384,-91,-126,-36,-139,-266,-168,-295,31,-134,-407,-95,-164,-151,-173,-330,-213,-259,86,-175,-461,-56,-127,-61,-180,-218,-177,-204,115,-165,-362,17,-129,-45,-57,-130,-80,-149,233,-1,-214,106,22,46,122,37,93,15,359,117,-118,280,170,198,216,116,134,124,407,221,-29,317,200,241,206,169,150,90,436,199,-55,285,208,272,200,98,116,26,318,100,-83,204,98,85,58,-11,25,-101,236,-3,-230,79,-31,27,-81,-167,-83,-228,187,-110,-428,-44,-123,-99,-182,-193,-188,-282,82,-203,-512,-76,-143,-147,-197,-257,-242,-279,37,-186,-453,13,-145,-134,-182,-175,-165,-226,109,-91,-364,-23,-87,12,-87,-129,-66,-98,282,-17,-240,107,73,164,20,52,64,5,381,155,-137,250,188,216,151,89,149,35,477,208,-85,303,183,237,190,168,206,66,493,221,-37,270,231,229,178,109,114,19,380,169,-156,176,112,119,71,-71,31,-65,296,56,-255,107,-46,-3,-75,-87,-98,-210,127,-134,-391,-56,-76,-111,-161,-215,-218,-237,52,-192,-489,-166,-131,-129,-215,-188,-189,-300,38,-189,-463,-47,-236,-114,-151,-242,-145,-242,133,-135,-353,27,-39,-29,-57,-109,-50,-96,257,12,-253,94,20,146,63,-16,14,16,340,155,-101,253,145,228,147,100,146,103,454,175,-58,339,253,231,200,163,203,119,409,243,-93,288,203,200,140,77,211,88,367,169,-106,169,73,160,74,-52,-37,-66,252,-44,-301,76,36,28,-70,-114,-146,-186,126,-181,-416,-61,-58,-72,-148,-281,-218,-333,64,-147,-485,-122,-156,-127,-186,-298,-252,-283,90,-245,-424,-70,-177,-154,-148,-276,-185,-261,98,-115,-320,36,-27,-43,-60,-114,-64,-132,283,1,-238,169,47,102,9,-2,93,-19,412,173,-102,253,210,225,165,88,143,105,460,224,-64,317,219,246,218,108,166,70,446,171,-26,290,183,210,154,110,133,58,388,147,-154,192,145,129,43,-44,3,-75,211,29,-302,83,20,30,-83,-134,-142,-99,150,-166,-316,-57,-135,-144,-184,-248,-259,-305,121,-183,-490,-93,-197,-114,-214,-241,-201,-340,84,-192,-448,-57,-185,-157,-180,-269,-189,-251,133,-145,-379,10,-101,-6,-81,-98,11,-138,289,7,-244,101,102,110,58,50,82,-28,375,145,-122,244,180,185,179,125,134,115,485,202,-75,281,251,229,239,128,172,157,511,189,-17,318,157,249,169,124,152,70,378,117,-179,191,164,140,112,-32,38,-88,240,9,-317,44,-18,6,-48,-73,-84,-187,140,-106,-392,-15,-122,-94,-151,-234,-220,-276,32,-187,-455,-112,-208,-172,-205,-264,-225,-278,16,-208,-498,-68,-175,-120,-116,-204,-213,-253,63,-120,-367,46,-32,45,-83,-83,-63,-145,149,-41,-208,154,111,147,71,36,45,42,402,135,-176,257,185,228,178,119,165,97,441,234,-55,261,239,235,185,190,229,72,457,164,-37,350,262,253,159,58,155,35,336,165,-111,256,115,143,83,-34,19,-35,263,34,-281,48,7,44,-82,-114,-136,-183,201,-101,-375,-36,-93,-115,-186,-261,-201,-267,18,-185,-437,-139,-201,-156,-153,-295,-225,-275,90,-209,-418,-101,-161,-122,-160,-196,-117,-229,95,-113,-353,-25,-71,-63,-76,-114,8,-134,184,2
--);

-- in=1000, out=1000, seno freq 0,009 + ruído em freq 0.03 e 0,02
--constant NOISY_ARRAY: T_NOISY_INPUT := (
--	11,21,31,40,48,56,62,67,70,72,73,73,72,69,66,62,58,53,48,44,40,36,33,31,29,29,29,30,32,35,38,42,46,49,53,57,59,62,63,64,63,62,59,56,51,46,40,33,26,19,11,4,-3,-10,-15,-21,-25,-28,-31,-32,-33,-33,-32,-30,-29,-26,-24,-22,-20,-19,-18,-18,-19,-21,-24,-27,-31,-37,-42,-49,-55,-62,-69,-75,-81,-86,-90,-93,-95,-96,-96,-93,-90,-85,-79,-72,-64,-55,-45,-35,-25,-16,-6,3,11,18,25,30,34,36,38,38,38,36,34,31,28,25,21,18,16,14,13,12,12,14,16,19,23,28,33,39,45,51,57,62,67,71,75,77,79,79,79,77,74,70,66,61,55,49,43,36,30,25,20,15,11,8,6,5,4,5,5,6,8,9,11,12,13,14,13,12,10,7,3,-2,-8,-15,-23,-31,-39,-48,-56,-65,-73,-80,-86,-92,-96,-99,-100,-100,-99,-96,-92,-87,-80,-73,-65,-57,-49,-41,-33,-25,-18,-12,-7,-3,-0,2,3,2,1,-1,-3,-6,-9,-12,-16,-18,-20,-22,-22,-22,-21,-18,-15,-11,-5,1,8,15,22,30,38,45,52,58,64,68,72,74,76,76,75,74,71,68,64,60,56,52,48,44,41,38,36,34,34,34,34,36,38,40,42,44,47,48,50,50,50,49,47,44,40,34,28,20,12,3,-6,-16,-26,-35,-45,-53,-61,-68,-74,-79,-82,-84,-84,-83,-81,-78,-74,-69,-63,-57,-51,-45,-39,-34,-29,-25,-22,-19,-18,-18,-19,-21,-24,-27,-31,-35,-40,-44,-48,-52,-55,-57,-58,-58,-58,-55,-52,-48,-42,-36,-29,-21,-13,-5,4,12,20,27,34,39,44,48,51,53,54,54,54,53,51,49,47,44,42,41,39,39,39,39,41,43,46,49,53,57,61,65,69,73,75,78,79,79,78,76,73,68,63,56,48,40,31,21,11,2,-8,-17,-25,-32,-39,-44,-48,-51,-52,-53,-52,-50,-47,-44,-40,-35,-31,-27,-23,-19,-16,-14,-13,-13,-14,-16,-19,-23,-28,-33,-39,-46,-52,-58,-64,-70,-75,-79,-82,-83,-84,-83,-81,-78,-74,-69,-63,-56,-48,-41,-33,-25,-17,-10,-4,2,7,12,15,18,19,20,20,20,20,19,18,17,16,16,17,18,19,22,25,29,34,39,45,51,57,64,70,75,80,85,88,90,91,91,90,87,83,78,72,65,58,50,41,33,24,17,9,3,-3,-8,-11,-14,-15,-15,-15,-13,-10,-7,-4,-0,4,7,10,13,15,15,15,14,11,8,3,-3,-9,-17,-24,-33,-41,-50,-58,-65,-72,-78,-83,-87,-90,-91,-91,-90,-88,-85,-80,-75,-70,-64,-57,-51,-45,-39,-34,-29,-25,-22,-19,-18,-17,-16,-16,-17,-18,-19,-20,-20,-20,-20,-19,-18,-15,-12,-7,-2,4,10,17,25,33,41,48,56,63,69,74,78,81,83,84,83,82,79,75,70,64,58,52,46,39,33,28,23,19,16,14,13,13,14,16,19,23,27,31,35,40,44,47,50,52,53,52,51,48,44,39,32,25,17,8,-2,-11,-21,-31,-40,-48,-56,-63,-68,-73,-76,-78,-79,-79,-78,-75,-73,-69,-65,-61,-57,-53,-49,-46,-43,-41,-39,-39,-39,-39,-41,-42,-44,-47,-49,-51,-53,-54,-54,-54,-53,-51,-48,-44,-39,-34,-27,-20,-12,-4,5,13,21,29,36,42,48,52,55,58,58,58,57,55,52,48,44,40,35,31,27,24,21,19,18,18,19,22,25,29,34,39,45,51,57,63,69,74,78,81,83,84,84,82,79,74,68,61,53,45,35,26,16,6,-3,-12,-20,-28,-34,-40,-44,-47,-49,-50,-50,-50,-48,-47,-44,-42,-40,-38,-36,-34,-34,-34,-34,-36,-38,-41,-44,-48,-52,-56,-60,-64,-68,-71,-74,-75,-76,-76,-74,-72,-68,-64,-58,-52,-45,-38,-30,-22,-15,-8,-1,5,11,15,18,21,22,22,22,20,18,16,12,9,6,3,1,-1,-2,-3,-2,0,3,7,12,18,25,33,41,49,57,65,73,80,87,92,96,99,100,100,99,96,92,86,80,73,65,56,48,39,31,23,15,8,2,-3,-7,-10,-12,-13,-14,-13,-12,-11,-9,-8,-6,-5,-5,-4,-5,-6,-8,-11,-15,-20,-25,-30,-36,-43,-49,-55,-61,-66,-70,-74,-77,-79,-79,-79,-77,-75,-71,-67,-62,-57,-51,-45,-39,-33,-28,-23,-19,-16,-14,-12,-12,-13,-14,-16,-18,-21,-25,-28,-31,-34,-36,-38,-38,-38,-36,-34,-30,-25,-18,-11,-3,6,16,25,35,45,55,64,72,79,85,90,93,96,96,95,93,90,86,81,75,69,62,55,49,42,37,31,27,24,21,19,18,18,19,20,22,24,26,29,30,32,33,33,32,31,28,25,21,15,10,3,-4,-11,-19,-26,-33,-40,-46,-51,-56,-59,-62,-63,-64,-63,-62,-59,-57,-53,-49,-46,-42,-38,-35,-32,-30,-29,-29,-29,-31,-33,-36,-40,-44,-48,-53,-58,-62,-66,-69,-72,-73,-73,-72,-70,-67,-62,-56,-48,-40,-31,-21,-11,-0
--);
	
-- L=64 cancelamento de ruído, funciona!
--constant COEFF_ARRAY : T_COEFF_INPUT := (
--	1,1,-1,-4,-8,-14,-18,-20,-21,-21,-20,-18,-15,-11,-7,-4,-1,2,4,4,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
--);
	
	component fir_filter 
	generic( 
		Win 		: INTEGER	; -- Input bit width
		Wmult 		: INTEGER	;-- Multiplier bit width 2*W1
		Wadd 		: INTEGER	;-- Adder width = Wmult+log2(L)-1
		Wout 		: INTEGER	;-- Output bit width
		BUTTON_HIGH : STD_LOGIC ;
		LFilter  	: INTEGER	);--Filter Length
	port (
		clk      : in  std_logic	;
		reset    : in  std_logic	;
		i_coeff  : in  ARRAY_COEFF(0 to Lfilter-1)		;
		i_data   : in  std_logic_vector( Win-1 	downto 0)	;
		o_data   : out std_logic_vector( Wout-1 downto 0)   ;
		read_out   : out integer  );
	end component;

	signal i_coeff 	: ARRAY_COEFF(0 to Lfilter-1); 
	signal i_data   : std_logic_vector( Win-1  downto 0);
	signal NOISY	: ARRAY_COEFF(0 to noisy_size-1);

begin
	
	u_fir_filter : fir_filter
	generic map( 
		Win 		 => Win				, -- Input bit width
		Wmult		 => Wmult			,
		Wadd		 => Wadd			,
		Wout 		 => Wout			,-- Output bit width
		BUTTON_HIGH  => BUTTON_HIGH		,
		LFilter  	 => LFilter			) -- Filter length	
	port map(
		clk         => clk       	,
		reset       => reset      	,
		i_coeff     => i_coeff		,
		i_data      => i_data 		,
		o_data     	=> o_data_buffer ,
		read_out  	=> read_out      );

	p_input : process (reset,clk)
		variable control  	: unsigned(11 downto 0):= (others=>'0');
		variable count 		: integer := 0;
		variable count2     : integer := 0;
		variable s			: integer RANGE 0 TO 2**8-1 :=255;
		variable first_time : std_logic := '0';
	begin
		if(reset=BUTTON_HIGH) then
			i_data       <= (others=>'0'); 
			count 		:= 0;
			count2 		:= 0;
			first_time	:='0';
			o_fir_coeff <= (others=>'0'); 
			o_input <= (others=>'0'); 
		elsif(rising_edge(clk)) then
			if(first_time='0') then
				for k in 0 to Lfilter-1 loop
					i_coeff(k)  <=  std_logic_vector(to_signed(COEFF_ARRAY(k),Win));
				end loop;			
				for j in 0 to noisy_size-1 loop
					NOISY(j)  <=  std_logic_vector(to_signed(NOISY_ARRAY(j),Win));
				end loop;
				first_time := '1';
			else
				--if(count>=5000 and count<10000) then
				--	s:= 0;
				--elsif (count>=10000) then 
				--	count:=0;
				--	s:=255;
				--end if;
				--i_data<=std_logic_vector(to_unsigned(s,Win));

				--count := count+1;
				--
				--if(count < 5000) then
				--	i_data   <= ('0',others=>'1');
				--elsif(count >= 5000 and count <10000) then
				--	i_data   <= (others=>'0');
				--elsif(count >=10000) then
				--	i_data   <= (others=>'0');
				--	count := 0;
				--end if;				
				--
				-- DELTA, STEP ...........
				--if(control=100 and count2 = 0) then  -- delta
				--	i_data       <= ('0',others=>'1');
				--elsif(control(11)='1' and count2 <3000 ) then  -- step
				--	i_data       <= ('0',others=>'1');
				--	count2 := count2 + 1;
				--else
				--	i_data       <= (others=>'0');
				--end if;
				--control := control + 1;
				------------------------------------------------

				-- DELTA, STEP, STEP, STEP, .......
				--if(control=10) then  -- delta
				--	i_data       <= ('0',others=>'1');
				--elsif(control(7)='1') then  -- step
				--	i_data       <= ('0',others=>'1');
				--else
				--	i_data       <= (others=>'0');
				--end if;
				--control := control + 1;
				-------------------------------------------------
				
				-- NOISY ANALOG SIGNAL
				if(count < noisy_size) then
					i_data <= NOISY(count);
					o_input <= NOISY(count);
					count := count + 1;
				else
					i_data <= (others=>'0');
				end if;
				-------------------------------------------------

				-- COEFFICIENTS
				if(count < Lfilter-1) then
					o_fir_coeff <= i_coeff(count);
				else
					o_fir_coeff <= (others=>'0');
				end if;
				---------------------------------------------------

				--count := count+1;
			end if;
		end if;
	end process p_input;
end rtl;
