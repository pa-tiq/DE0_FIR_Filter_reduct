LIBRARY work;
USE work.n_bit_int.ALL;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fir_filter_test is
	generic( 
		Win 			: INTEGER 	; -- Input bit width
		Wmult			: INTEGER 	;-- Multiplier bit width 2*W1
		Wadd 			: INTEGER 	;-- Adder width = Wmult+log2(L)-1
		Wout 			: INTEGER 	;-- Output bit width
		BUTTON_HIGH 	: STD_LOGIC ;
		PATTERN_SIZE	: INTEGER 	;
		RANGE_LOW 		: INTEGER 	; --pattern range: power of 2
		RANGE_HIGH 		: INTEGER 	; --must change pattern too
		LFilter  		: INTEGER 	); -- Filter length
	port (
		clk              	  : in  std_logic;
		reset                 : in  std_logic;
		o_data_buffer         : out std_logic_vector( Wout-1 downto 0);
		o_fir_coeff           : out std_logic_vector( Win-1 downto 0);
		read_out              : out integer );
end fir_filter_test;

architecture rtl of fir_filter_test is

	constant noisy_size : integer := 1060;
	type T_NOISY_INPUT is array(0 to noisy_size-1) of integer range RANGE_LOW to RANGE_HIGH;
	type T_COEFF_INPUT is array(0 to LFilter-1) of integer range RANGE_LOW to RANGE_HIGH;

	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--0,1,2,5,9,16,25,36,48,62,77,92,105,115,123,127,127,123,115,
	--105,92,77,62,48,36,25,16,9,5,2,1,0);

	-- L=256 RANGE -256 TO 255
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,-1,-1,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,
	--	-2,-2,-1,0,1,2,3,4,5,6,7,8,10,11,12,13,14,15,15,16,17,17,17,17,17,16,16,15,14,12,
	--	11,9,7,5,3,0,-3,-6,-9,-12,-15,-18,-21,-24,-27,-30,-33,-35,-38,-40,-42,-43,-45,-45,
	--	-46,-45,-45,-44,-42,-39,-37,-33,-29,-24,-19,-13,-7,0,8,16,24,33,42,52,62,73,83,94,
	--	105,116,127,137,148,159,169,179,188,197,206,214,221,228,234,240,244,248,251,253,255,
	--	255,253,251,248,244,240,234,228,221,214,206,197,188,179,169,159,148,137,127,116,105,
	--	94,83,73,62,52,42,33,24,16,8,0,-7,-13,-19,-24,-29,-33,-37,-39,-42,-44,-45,-45,-46,-45,
	--	-45,-43,-42,-40,-38,-35,-33,-30,-27,-24,-21,-18,-15,-12,-9,-6,-3,0,3,5,7,9,11,12,14,
	--	15,16,16,17,17,17,17,17,16,15,15,14,13,12,11,10,8,7,6,5,4,3,2,1,0,-1,-2,-2,-3,-3,-4,
	--	-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,-1,-1,0,0,0,0,0,0);

	-- L=256 RANGE -512 TO 511
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,-1,-1,-2,-2,-3,-4,-4,-5,-5,-6,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-7,-6,-5,-4,-3,
	--	-2,0,2,4,6,8,10,12,15,17,19,22,24,26,28,29,31,32,33,34,34,34,34,33,31,30,27,25,22,18,14,
	--	10,5,0,-5,-11,-17,-23,-29,-36,-42,-48,-54,-60,-66,-71,-76,-80,-84,-87,-89,-91,-91,-91,
	--	-90,-87,-84,-79,-74,-67,-58,-49,-39,-27,-14,0,15,31,48,66,85,105,125,146,167,189,210,232,
	--	254,276,298,319,339,359,378,396,414,430,445,459,471,482,491,498,504,509,511,511,509,504,
	--	498,491,482,471,459,445,430,414,396,378,359,339,319,298,276,254,232,210,189,167,146,125,
	--	105,85,66,48,31,15,0,-14,-27,-39,-49,-58,-67,-74,-79,-84,-87,-90,-91,-91,-91,-89,-87,-84,
	--	-80,-76,-71,-66,-60,-54,-48,-42,-36,-29,-23,-17,-11,-5,0,5,10,14,18,22,25,27,30,31,33,34,
	--	34,34,34,33,32,31,29,28,26,24,22,19,17,15,12,10,8,6,4,2,0,-2,-3,-4,-5,-6,-7,-8,-8,-8,-8,
	--	-8,-8,-8,-8,-7,-7,-6,-5,-5,-4,-4,-3,-2,-2,-1,-1,-1,0,0,0,0,0);

	-- L=256 RANGE -512 TO 511
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,1,0,-1,0,1,1,0,-1,-1,1,1,0,-1,-1,1,1,0,-1,-1,1,
	--	2,0,-2,-1,1,2,0,-2,-1,1,3,0,-3,-2,2,3,0,-3,-2,2,4,0,-4,-3,3,4,0,-5,-3,3,5,0,-6,-4,4,6,0,-7,-4,4,7,0,
	--	-8,-5,5,9,0,-10,-6,6,11,0,-12,-8,8,14,0,-15,-10,10,17,0,-19,-13,14,23,0,-27,-18,20,35,0,-43,-30,34,
	--	64,0,-97,-80,119,387,511,511,387,119,-80,-97,0,64,34,-30,-43,0,35,20,-18,-27,0,23,14,-13,-19,0,17,10,
	--	-10,-15,0,14,8,-8,-12,0,11,6,-6,-10,0,9,5,-5,-8,0,7,4,-4,-7,0,6,4,-4,-6,0,5,3,-3,-5,0,4,3,-3,-4,0,4,2,
	--	-2,-3,0,3,2,-2,-3,0,3,1,-1,-2,0,2,1,-1,-2,0,2,1,-1,-1,0,1,1,-1,-1,0,1,1,-1,-1,0,1,1,0,-1,0,1,0,0,-1,0,
	--	1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
	
	-- L=512 RANGE 256 TO 255
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-3,
	--	-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,
	--	-4,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,0,0,0,1,1,2,2,3,3,4,4,5,6,6,7,7,8,8,9,10,
	--	10,11,11,12,12,13,13,14,14,15,15,15,16,16,16,17,17,17,17,17,17,17,17,17,17,
	--	16,16,16,15,15,14,14,13,12,12,11,10,9,8,7,6,5,4,3,1,0,-1,-3,-4,-6,-7,-9,-10,
	--	-12,-13,-15,-16,-18,-19,-21,-23,-24,-26,-27,-29,-30,-31,-33,-34,-35,-37,-38,
	--	-39,-40,-41,-42,-43,-43,-44,-45,-45,-45,-45,-46,-46,-45,-45,-45,-44,-44,-43,
	--	-42,-41,-40,-38,-37,-35,-33,-31,-29,-27,-24,-22,-19,-16,-13,-10,-7,-4,0,4,8,
	--	11,16,20,24,28,33,38,42,47,52,57,62,67,73,78,83,89,94,99,105,110,116,121,127,
	--	132,137,143,148,153,159,164,169,174,179,184,188,193,197,202,206,210,214,218,
	--	222,225,228,231,234,237,240,242,244,246,248,250,251,252,253,254,255,255,255,
	--	255,254,253,252,251,250,248,246,244,242,240,237,234,231,228,225,222,218,214,
	--	210,206,202,197,193,188,184,179,174,169,164,159,153,148,143,137,132,127,121,
	--	116,110,105,99,94,89,83,78,73,67,62,57,52,47,42,38,33,28,24,20,16,11,8,4,0,
	--	-4,-7,-10,-13,-16,-19,-22,-24,-27,-29,-31,-33,-35,-37,-38,-40,-41,-42,-43,-44,
	--	-44,-45,-45,-45,-46,-46,-45,-45,-45,-45,-44,-43,-43,-42,-41,-40,-39,-38,-37,
	--	-35,-34,-33,-31,-30,-29,-27,-26,-24,-23,-21,-19,-18,-16,-15,-13,-12,-10,-9,-7,
	--	-6,-4,-3,-1,0,1,3,4,5,6,7,8,9,10,11,12,12,13,14,14,15,15,16,16,16,17,17,17,17,
	--	17,17,17,17,17,17,16,16,16,15,15,15,14,14,13,13,12,12,11,11,10,10,9,8,8,7,7,6,
	--	6,5,4,4,3,3,2,2,1,1,0,0,0,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,
	--	-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-1,-1,
	--	-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0);

	-- L=512 RANGE -512 TO 511 (1)
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,0,0,-1,-1,-1,-2,-2,-1,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,0,1,1,2,3,3,3,2,1,0,-1,-2,-3,-3,-3,-3,-3,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-4,-5,-5,-5,-4,-3,-1,1,2,4,5,6,6,5,3,2,-1,-3,-5,-6,-7,-7,-6,-4,-2,0,3,5,7,8,8,7,5,3,0,-3,-6,-8,-9,-9,-8,-6,-3,0,4,7,9,11,11,10,8,4,0,-4,-8,-11,-13,-13,-12,-9,-6,-1,4,9,12,15,15,14,11,7,2,-4,-10,-14,-17,-18,-17,-14,-9,-3,4,11,17,21,22,21,17,11,4,-5,-13,-20,-25,-27,-26,-22,-15,-6,5,15,24,31,34,33,28,20,8,-5,-18,-30,-40,-45,-44,-39,-28,-13,5,24,41,55,63,64,57,43,21,-5,-34,-63,-87,-104,-110,-104,-82,-46,5,68,139,216,292,363,424,471,501,511,511,501,471,424,363,292,216,139,68,5,-46,-82,-104,-110,-104,-87,-63,-34,-5,21,43,57,64,63,55,41,24,5,-13,-28,-39,-44,-45,-40,-30,-18,-5,8,20,28,33,34,31,24,15,5,-6,-15,-22,-26,-27,-25,-20,-13,-5,4,11,17,21,22,21,17,11,4,-3,-9,-14,-17,-18,-17,-14,-10,-4,2,7,11,14,15,15,12,9,4,-1,-6,-9,-12,-13,-13,-11,-8,-4,0,4,8,10,11,11,9,7,4,0,-3,-6,-8,-9,-9,-8,-6,-3,0,3,5,7,8,8,7,5,3,0,-2,-4,-6,-7,-7,-6,-5,-3,-1,2,3,5,6,6,5,4,2,1,-1,-3,-4,-5,-5,-5,-4,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-3,-3,-3,-3,-3,-2,-1,0,1,2,3,3,3,2,1,1,0,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-1,-2,-2,-1,-1,-1,0,0,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,-1,0,0,0,0,0
	--);
	
    -- L=512 RANGE -512 TO 511 SEM JANELA
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	4,3,1,-1,-3,-4,-4,-4,-3,-1,1,3,4,4,4,2,0,-2,-4,-5,-4,-3,-1,1,3,4,5,4,3,1,-1,-3,-5,-5,-4,-2,0,2,4,5,5,4,2,-1,-3,-5,-5,-5,-3,-1,2,4,5,5,4,2,0,-2,-4,-5,-5,-4,-2,1,3,5,6,5,3,1,-2,-4,-6,-6,-5,-3,0,3,5,6,6,4,2,-1,-4,-6,-6,-6,-4,-1,2,5,6,7,5,3,0,-3,-6,-7,-7,-5,-2,1,4,6,7,6,4,1,-2,-5,-7,-7,-6,-3,0,4,6,8,8,6,3,-1,-5,-7,-8,-7,-5,-1,3,6,8,9,7,4,0,-4,-7,-9,-9,-7,-3,2,6,9,10,9,6,2,-3,-7,-10,-10,-9,-5,0,5,9,11,11,8,4,-2,-7,-11,-12,-11,-7,-2,4,9,12,13,11,6,0,-6,-11,-14,-14,-10,-5,2,9,14,15,14,9,3,-5,-12,-16,-17,-14,-8,0,8,15,19,18,14,6,-3,-12,-19,-22,-20,-13,-4,7,17,23,25,21,12,0,-13,-23,-29,-29,-22,-10,5,20,31,36,33,23,6,-13,-31,-43,-47,-40,-23,0,26,49,63,64,51,24,-13,-53,-88,-108,-107,-80,-24,56,153,258,357,439,492,511,492,439,357,258,153,56,-24,-80,-107,-108,-88,-53,-13,24,51,64,63,49,26,0,-23,-40,-47,-43,-31,-13,6,23,33,36,31,20,5,-10,-22,-29,-29,-23,-13,0,12,21,25,23,17,7,-4,-13,-20,-22,-19,-12,-3,6,14,18,19,15,8,0,-8,-14,-17,-16,-12,-5,3,9,14,15,14,9,2,-5,-10,-14,-14,-11,-6,0,6,11,13,12,9,4,-2,-7,-11,-12,-11,-7,-2,4,8,11,11,9,5,0,-5,-9,-10,-10,-7,-3,2,6,9,10,9,6,2,-3,-7,-9,-9,-7,-4,0,4,7,9,8,6,3,-1,-5,-7,-8,-7,-5,-1,3,6,8,8,6,4,0,-3,-6,-7,-7,-5,-2,1,4,6,7,6,4,1,-2,-5,-7,-7,-6,-3,0,3,5,7,6,5,2,-1,-4,-6,-6,-6,-4,-1,2,4,6,6,5,3,0,-3,-5,-6,-6,-4,-2,1,3,5,6,5,3,1,-2,-4,-5,-5,-4,-2,0,2,4,5,5,4,2,-1,-3,-5,-5,-5,-3,-1,2,4,5,5,4,2,0,-2,-4,-5,-5,-3,-1,1,3,4,5,4,3,1,-1,-3,-4,-5,-4,-2,0,2,4,4,4,3,1,-1,-3,-4,-4,-4,-3,-1,1,3
	--);	
	
	-- L=512 RANGE -512 TO 511 (hamming) b=0.15
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,0,0,-1,-1,-1,-2,-2,-1,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,0,1,1,2,3,3,3,2,1,0,-1,-2,-3,-3,-3,-3,-3,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-4,-5,-5,-5,-4,-3,-1,1,2,4,5,6,6,5,3,2,-1,-3,-5,-6,-7,-7,-6,-4,-2,0,3,5,7,8,8,7,5,3,0,-3,-6,-8,-9,-9,-8,-6,-3,0,4,7,9,11,11,10,8,4,0,-4,-8,-11,-13,-13,-12,-9,-6,-1,4,9,12,15,15,14,11,7,2,-4,-10,-14,-17,-18,-17,-14,-9,-3,4,11,17,21,22,21,17,11,4,-5,-13,-20,-25,-27,-26,-22,-15,-6,5,15,24,31,34,33,28,20,8,-5,-18,-30,-40,-45,-44,-39,-28,-13,5,24,41,55,63,64,57,43,21,-5,-34,-63,-87,-104,-110,-104,-82,-46,5,68,139,216,292,363,424,471,501,511,511,501,471,424,363,292,216,139,68,5,-46,-82,-104,-110,-104,-87,-63,-34,-5,21,43,57,64,63,55,41,24,5,-13,-28,-39,-44,-45,-40,-30,-18,-5,8,20,28,33,34,31,24,15,5,-6,-15,-22,-26,-27,-25,-20,-13,-5,4,11,17,21,22,21,17,11,4,-3,-9,-14,-17,-18,-17,-14,-10,-4,2,7,11,14,15,15,12,9,4,-1,-6,-9,-12,-13,-13,-11,-8,-4,0,4,8,10,11,11,9,7,4,0,-3,-6,-8,-9,-9,-8,-6,-3,0,3,5,7,8,8,7,5,3,0,-2,-4,-6,-7,-7,-6,-5,-3,-1,2,3,5,6,6,5,4,2,1,-1,-3,-4,-5,-5,-5,-4,-2,-1,1,2,3,4,4,4,3,2,1,-1,-2,-3,-3,-3,-3,-3,-2,-1,0,1,2,3,3,3,2,1,1,0,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,2,2,2,1,1,0,-1,-1,-1,-2,-2,-1,-1,-1,0,0,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,-1,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (hamming) b=0.05
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,1,1,1,0,0,-1,-1,-2,-2,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-2,-2,-1,0,0,1,2,3,3,4,5,5,5,6,6,6,5,5,4,4,3,2,1,0,-2,-3,-4,-5,-6,-7,-8,-9,-9,-9,-9,-9,-9,-8,-7,-6,-5,-4,-2,0,1,3,5,7,8,10,11,12,12,13,13,13,12,11,10,8,6,4,2,0,-3,-5,-8,-10,-13,-15,-16,-18,-19,-19,-19,-19,-18,-17,-15,-13,-10,-7,-4,0,3,7,10,14,17,20,22,24,26,27,27,26,25,23,21,17,14,9,5,0,-6,-11,-16,-21,-25,-30,-33,-36,-38,-39,-40,-39,-37,-35,-31,-26,-21,-15,-8,0,7,15,23,30,37,44,49,54,57,59,60,59,57,53,47,40,32,22,11,0,-13,-26,-38,-51,-63,-75,-85,-94,-101,-106,-108,-108,-105,-99,-90,-79,-63,-45,-24,0,26,55,86,118,152,187,221,256,291,324,356,386,413,438,460,478,492,503,509,511,511,509,503,492,478,460,438,413,386,356,324,291,256,221,187,152,118,86,55,26,0,-24,-45,-63,-79,-90,-99,-105,-108,-108,-106,-101,-94,-85,-75,-63,-51,-38,-26,-13,0,11,22,32,40,47,53,57,59,60,59,57,54,49,44,37,30,23,15,7,0,-8,-15,-21,-26,-31,-35,-37,-39,-40,-39,-38,-36,-33,-30,-25,-21,-16,-11,-6,0,5,9,14,17,21,23,25,26,27,27,26,24,22,20,17,14,10,7,3,0,-4,-7,-10,-13,-15,-17,-18,-19,-19,-19,-19,-18,-16,-15,-13,-10,-8,-5,-3,0,2,4,6,8,10,11,12,13,13,13,12,12,11,10,8,7,5,3,1,0,-2,-4,-5,-6,-7,-8,-9,-9,-9,-9,-9,-9,-8,-7,-6,-5,-4,-3,-2,0,1,2,3,4,4,5,5,6,6,6,5,5,5,4,3,3,2,1,0,0,-1,-2,-2,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-2,-2,-1,-1,0,0,1,1,1,2,2,2,2,2,2,2,2,2,1,1,1,1,0,0,0,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0
	--);
	
	-- L=512 RANGE -512 TO 511 (hamming) b=0.01
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-5,-5,-6,-6,-7,-7,-8,-9,-9,-10,-11,-11,-12,-13,-14,-14,-15,-16,-17,-18,-19,-20,-21,-22,-23,-24,-25,-26,-27,-28,-29,-30,-31,-32,-33,-34,-35,-37,-38,-39,-40,-41,-42,-43,-44,-45,-46,-47,-48,-49,-50,-51,-52,-53,-54,-54,-55,-56,-57,-57,-58,-58,-59,-59,-59,-60,-60,-60,-60,-60,-60,-59,-59,-59,-58,-58,-57,-56,-56,-55,-54,-52,-51,-50,-48,-47,-45,-43,-41,-39,-37,-35,-33,-30,-27,-25,-22,-19,-16,-12,-9,-5,-2,2,6,10,14,18,23,27,32,37,42,47,52,57,62,68,73,79,85,91,97,103,109,115,121,128,134,141,148,154,161,168,175,182,189,196,203,210,217,224,231,238,246,253,260,267,274,282,289,296,303,310,317,324,331,338,344,351,358,364,371,377,383,390,396,402,407,413,419,424,430,435,440,445,450,454,459,463,467,471,475,478,482,485,488,491,494,496,499,501,503,504,506,507,508,509,510,511,511,511,511,510,509,508,507,506,504,503,501,499,496,494,491,488,485,482,478,475,471,467,463,459,454,450,445,440,435,430,424,419,413,407,402,396,390,383,377,371,364,358,351,344,338,331,324,317,310,303,296,289,282,274,267,260,253,246,238,231,224,217,210,203,196,189,182,175,168,161,154,148,141,134,128,121,115,109,103,97,91,85,79,73,68,62,57,52,47,42,37,32,27,23,18,14,10,6,2,-2,-5,-9,-12,-16,-19,-22,-25,-27,-30,-33,-35,-37,-39,-41,-43,-45,-47,-48,-50,-51,-52,-54,-55,-56,-56,-57,-58,-58,-59,-59,-59,-60,-60,-60,-60,-60,-60,-59,-59,-59,-58,-58,-57,-57,-56,-55,-54,-54,-53,-52,-51,-50,-49,-48,-47,-46,-45,-44,-43,-42,-41,-40,-39,-38,-37,-35,-34,-33,-32,-31,-30,-29,-28,-27,-26,-25,-24,-23,-22,-21,-20,-19,-18,-17,-16,-15,-14,-14,-13,-12,-11,-11,-10,-9,-9,-8,-7,-7,-6,-6,-5,-5,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.1
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,1,1,1,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,2,3,3,3,2,2,1,0,-1,-2,-3,-3,-4,-4,-3,-2,-1,0,1,3,4,4,5,5,4,3,2,0,-2,-3,-5,-6,-6,-6,-5,-4,-2,0,2,4,6,7,8,7,6,5,3,0,-3,-5,-7,-9,-10,-9,-8,-6,-3,0,3,7,9,11,12,12,10,8,4,0,-4,-8,-12,-14,-15,-15,-13,-10,-5,0,5,11,15,18,19,19,16,12,7,0,-7,-13,-19,-23,-24,-24,-21,-16,-8,0,9,17,24,29,32,31,27,20,11,0,-12,-23,-33,-40,-43,-42,-37,-28,-15,0,16,33,47,57,63,62,55,42,23,0,-26,-52,-76,-95,-107,-109,-100,-79,-45,0,56,119,187,257,325,386,438,478,503,511,511,503,478,438,386,325,257,187,119,56,0,-45,-79,-100,-109,-107,-95,-76,-52,-26,0,23,42,55,62,63,57,47,33,16,0,-15,-28,-37,-42,-43,-40,-33,-23,-12,0,11,20,27,31,32,29,24,17,9,0,-8,-16,-21,-24,-24,-23,-19,-13,-7,0,7,12,16,19,19,18,15,11,5,0,-5,-10,-13,-15,-15,-14,-12,-8,-4,0,4,8,10,12,12,11,9,7,3,0,-3,-6,-8,-9,-10,-9,-7,-5,-3,0,3,5,6,7,8,7,6,4,2,0,-2,-4,-5,-6,-6,-6,-5,-3,-2,0,2,3,4,5,5,4,4,3,1,0,-1,-2,-3,-4,-4,-3,-3,-2,-1,0,1,2,2,3,3,3,2,1,1,0,-1,-1,-2,-2,-2,-2,-2,-1,-1,0,1,1,1,1,1,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	
	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.05
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,1,1,1,2,2,2,2,2,3,3,3,2,2,2,2,1,1,1,0,-1,-1,-2,-2,-3,-3,-4,-4,-5,-5,-5,-5,-5,-4,-4,-3,-3,-2,-1,0,1,2,3,4,5,6,7,7,8,8,8,8,8,7,7,6,4,3,2,0,-2,-3,-5,-7,-8,-10,-11,-12,-13,-14,-14,-13,-13,-12,-11,-9,-7,-5,-3,0,3,6,8,11,14,16,18,20,21,22,22,21,21,19,17,15,12,8,4,0,-4,-9,-13,-17,-22,-25,-28,-31,-33,-34,-35,-34,-33,-30,-27,-23,-18,-13,-7,0,7,14,21,28,35,41,46,50,54,56,56,56,54,50,45,39,31,21,11,0,-12,-24,-37,-49,-61,-72,-82,-91,-98,-103,-105,-105,-103,-97,-89,-77,-62,-44,-24,0,26,55,85,118,151,186,221,256,290,323,355,385,413,438,459,478,492,503,509,511,511,509,503,492,478,459,438,413,385,355,323,290,256,221,186,151,118,85,55,26,0,-24,-44,-62,-77,-89,-97,-103,-105,-105,-103,-98,-91,-82,-72,-61,-49,-37,-24,-12,0,11,21,31,39,45,50,54,56,56,56,54,50,46,41,35,28,21,14,7,0,-7,-13,-18,-23,-27,-30,-33,-34,-35,-34,-33,-31,-28,-25,-22,-17,-13,-9,-4,0,4,8,12,15,17,19,21,21,22,22,21,20,18,16,14,11,8,6,3,0,-3,-5,-7,-9,-11,-12,-13,-13,-14,-14,-13,-12,-11,-10,-8,-7,-5,-3,-2,0,2,3,4,6,7,7,8,8,8,8,8,7,7,6,5,4,3,2,1,0,-1,-2,-3,-3,-4,-4,-5,-5,-5,-5,-5,-4,-4,-3,-3,-2,-2,-1,-1,0,1,1,1,2,2,2,2,3,3,3,2,2,2,2,2,1,1,1,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 (BLACKMAN) b=0.01
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-4,-4,-5,-5,-5,-6,-6,-7,-7,-8,-8,-9,-9,-10,-10,-11,-11,-12,-12,-13,-14,-14,-15,-16,-16,-17,-18,-18,-19,-20,-21,-21,-22,-23,-23,-24,-25,-25,-26,-27,-27,-28,-29,-29,-30,-30,-31,-31,-32,-32,-32,-33,-33,-33,-34,-34,-34,-34,-34,-34,-33,-33,-33,-33,-32,-32,-31,-30,-29,-29,-28,-27,-25,-24,-23,-21,-20,-18,-16,-14,-12,-10,-8,-6,-3,0,2,5,8,11,15,18,22,25,29,33,37,41,46,50,55,59,64,69,74,79,85,90,96,101,107,113,119,125,131,138,144,151,157,164,171,178,184,191,198,206,213,220,227,234,242,249,256,264,271,278,286,293,300,307,315,322,329,336,343,350,357,364,370,377,384,390,396,403,409,415,421,426,432,437,443,448,453,457,462,466,471,475,478,482,485,489,492,495,497,500,502,504,505,507,508,509,510,511,511,511,511,510,509,508,507,505,504,502,500,497,495,492,489,485,482,478,475,471,466,462,457,453,448,443,437,432,426,421,415,409,403,396,390,384,377,370,364,357,350,343,336,329,322,315,307,300,293,286,278,271,264,256,249,242,234,227,220,213,206,198,191,184,178,171,164,157,151,144,138,131,125,119,113,107,101,96,90,85,79,74,69,64,59,55,50,46,41,37,33,29,25,22,18,15,11,8,5,2,0,-3,-6,-8,-10,-12,-14,-16,-18,-20,-21,-23,-24,-25,-27,-28,-29,-29,-30,-31,-32,-32,-33,-33,-33,-33,-34,-34,-34,-34,-34,-34,-33,-33,-33,-32,-32,-32,-31,-31,-30,-30,-29,-29,-28,-27,-27,-26,-25,-25,-24,-23,-23,-22,-21,-21,-20,-19,-18,-18,-17,-16,-16,-15,-14,-14,-13,-12,-12,-11,-11,-10,-10,-9,-9,-8,-8,-7,-7,-6,-6,-5,-5,-5,-4,-4,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- L=512 RANGE -512 TO 511 ofdm
	constant COEFF_ARRAY : T_COEFF_INPUT := (
		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,-1,0,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-2,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-2,2,0,-3,1,2,-2,-1,3,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-4,1,3,-3,-2,4,-1,-4,3,2,-5,0,5,-3,-3,5,0,-5,3,4,-6,0,6,-3,-4,6,1,-7,3,6,-7,-2,8,-3,-7,8,3,-10,4,9,-9,-4,13,-4,-12,11,6,-17,4,17,-15,-10,24,-4,-27,23,20,-44,4,64,-56,-77,261,511,261,-77,-56,64,4,-44,20,23,-27,-4,24,-10,-15,17,4,-17,6,11,-12,-4,13,-4,-9,9,4,-10,3,8,-7,-3,8,-2,-7,6,3,-7,1,6,-4,-3,6,0,-6,4,3,-5,0,5,-3,-3,5,0,-5,2,3,-4,-1,4,-2,-3,3,1,-4,1,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,3,-1,-2,2,1,-3,0,2,-2,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,1,0,-2,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,0,-1,0,1,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	);

	-- L=2048 RANGE -127 to 126 HAMMING
	--constant COEFF_ARRAY : T_COEFF_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,4,4,4,4,4,4,4,3,3,3,3,3,3,2,2,2,2,2,1,1,1,1,1,0,0,0,0,0,-1,-1,-1,-1,-2,-2,-2,-2,-3,-3,-3,-3,-3,-4,-4,-4,-4,-5,-5,-5,-5,-5,-6,-6,-6,-6,-6,-7,-7,-7,-7,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-8,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-8,-8,-8,-8,-8,-8,-8,-8,-7,-7,-7,-7,-7,-6,-6,-6,-6,-5,-5,-5,-5,-4,-4,-4,-4,-3,-3,-3,-2,-2,-2,-1,-1,-1,0,0,0,1,1,1,2,2,2,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,11,12,12,12,12,12,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,13,13,13,13,13,12,12,12,12,11,11,11,10,10,10,9,9,9,8,8,7,7,6,6,5,5,4,4,3,3,2,2,1,1,0,-1,-1,-2,-2,-3,-4,-4,-5,-6,-6,-7,-7,-8,-9,-9,-10,-11,-11,-12,-12,-13,-14,-14,-15,-15,-16,-16,-17,-18,-18,-19,-19,-20,-20,-21,-21,-22,-22,-22,-23,-23,-24,-24,-24,-25,-25,-25,-25,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-25,-25,-25,-25,-24,-24,-24,-23,-23,-22,-22,-21,-21,-20,-19,-19,-18,-17,-16,-16,-15,-14,-13,-12,-11,-10,-9,-8,-7,-6,-5,-4,-2,-1,0,1,2,4,5,6,8,9,11,12,14,15,17,18,20,21,23,24,26,28,29,31,33,34,36,38,39,41,43,44,46,48,50,51,53,55,57,58,60,62,64,65,67,69,70,72,74,75,77,79,80,82,84,85,87,88,90,91,93,94,96,97,99,100,101,103,104,105,106,108,109,110,111,112,113,114,115,116,117,118,119,120,120,121,122,122,123,123,124,124,125,125,126,126,126,126,127,127,127,127,127,127,127,127,126,126,126,126,125,125,124,124,123,123,122,122,121,120,120,119,118,117,116,115,114,113,112,111,110,109,108,106,105,104,103,101,100,99,97,96,94,93,91,90,88,87,85,84,82,80,79,77,75,74,72,70,69,67,65,64,62,60,58,57,55,53,51,50,48,46,44,43,41,39,38,36,34,33,31,29,28,26,24,23,21,20,18,17,15,14,12,11,9,8,6,5,4,2,1,0,-1,-2,-4,-5,-6,-7,-8,-9,-10,-11,-12,-13,-14,-15,-16,-16,-17,-18,-19,-19,-20,-21,-21,-22,-22,-23,-23,-24,-24,-24,-25,-25,-25,-25,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-26,-25,-25,-25,-25,-24,-24,-24,-23,-23,-22,-22,-22,-21,-21,-20,-20,-19,-19,-18,-18,-17,-16,-16,-15,-15,-14,-14,-13,-12,-12,-11,-11,-10,-9,-9,-8,-7,-7,-6,-6,-5,-4,-4,-3,-2,-2,-1,-1,0,1,1,2,2,3,3,4,4,5,5,6,6,7,7,8,8,9,9,9,10,10,10,11,11,11,12,12,12,12,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,13,13,13,13,13,12,12,12,12,12,11,11,11,11,10,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,2,2,2,1,1,1,0,0,0,-1,-1,-1,-2,-2,-2,-3,-3,-3,-4,-4,-4,-4,-5,-5,-5,-5,-6,-6,-6,-6,-7,-7,-7,-7,-7,-8,-8,-8,-8,-8,-8,-8,-8,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-9,-8,-8,-8,-8,-8,-8,-8,-8,-8,-7,-7,-7,-7,-7,-7,-6,-6,-6,-6,-6,-5,-5,-5,-5,-5,-4,-4,-4,-4,-3,-3,-3,-3,-3,-2,-2,-2,-2,-1,-1,-1,-1,0,0,0,0,0,1,1,1,1,1,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,3,3,3,3,3,3,3,2,2,2,2,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-4,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-3,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- noisy sin -127 to 126
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-10,1,11,35,36,18,49,41,42,51,51,56,70,75,79,79,72,87,96,93,100,
	--	101,98,104,100,111,101,103,106,95,121,115,109,121,103,111,109,111,
	--	110,101,104,101,103,103,100,85,87,76,73,75,80,62,64,56,59,41,42,40,
	--	38,35,21,6,5,-3,11,-11,-9,-20,-19,-35,-44,-49,-43,-52,-58,-53,-64,
	--	-70,-66,-84,-80,-83,-93,-93,-105,-108,-103,-102,-94,-114,-111,-114,
	--	-126,-119,-127,-112,-122,-117,-120,-114);

	--noisy sawtooth -64 to 63
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-30,-25,-33,-32,-20,-46,-30,-35,-26,-15,-12,-27,-20,-13,-15,-8 ,-6 ,-16,-8 ,-24,7  ,-7 ,-11,0  ,-9 ,5  ,2  ,28 ,20 ,-11,17 ,2  ,14 ,19 ,26 ,19 ,37 ,20 ,29 ,33 ,30 ,39 ,35 ,27 ,19 ,54 ,33 ,41 ,47 ,44 ,37 ,42 ,47 ,63 ,44 ,60 ,57 ,54 ,48 ,57 ,60 ,50 ,-35,-42,-34,-29,-38,-31,-24,-42,-14,0  ,-12,-22,-13,-25,3  ,-4 ,-4 ,-17,-5 ,-11,-7 ,-8 ,-10,-8 ,0  ,-12,11 ,6  ,15 ,13 ,16 ,0  ,6  ,12 ,19 ,30 ,19 ,34
	--	);

	--noisy sawtooth -256 to 255
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-155,-124,-155,-177,-200,-134,-104,-138,-140,-125,-147,-119,-102,-87 ,-85 ,-54 ,-65 ,2   ,-45 ,15  ,-70 ,-18 ,-40 ,-3  ,3   ,-90 ,-53 ,-50 ,22  ,67  ,9   ,56  ,53  ,2   ,61  ,26  ,114 ,64  ,131 ,63  ,106 ,89  ,25  ,69  ,133 ,115 ,83  ,107 ,145 ,107 ,184 ,132 ,227 ,130 ,182 ,127 ,162 ,173 ,215 ,241 ,224 ,206 ,256 ,-142,-160,-138,-137,-181,-112,-156,-148,-113,-124,-112,-79 ,-56 ,-95 ,-69 ,-83 ,-60 ,-46 ,-78 ,-39 ,-21 ,-33 ,32  ,-45 ,-43 ,-73 ,29  ,34  ,6   ,48  ,28  ,39  ,39  ,57  ,51  ,154 ,18		
	--);

	-- TAMANHO 1060 - Símbolo OFDM parte real, -512 to 511
	constant NOISY_ARRAY : T_NOISY_INPUT := (
		49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,-8,-252,-50,257,131,-90,5,157,127,28,-93,-149,13,112,-163,-382,-122,189,158,75,50,-166,-386,-280,-62,56,178,156,-138,-239,35,83,-201,-143,231,201,-134,-148,1,-117,-248,-126,-9,2,87,129,-59,-271,-297,-202,-33,141,83,-163,-215,-66,-97,-263,-163,123,159,-20,-31,131,200,217,341,368,100,-137,-28,131,38,-18,179,270,60,-114,-110,-115,-81,52,-8,-247,-187,132,176,39,121,92,-338,-512,-44,336,189,63,176,112,-90,-67,20,-13,69,172,-87,-376,-133,229,58,-304,-288,-133,-161,-152,-17,-24,-148,-149,-103,-160,-203,-158,-129,-90,43,175,221,202,51,-220,-289,-14,210,91,-72,3,85,-48,-167,-25,196,187,-7,-75,77,226,197,58,-77,-135,-26,191,227,19,-99,13,48,-119,-185,-14,138,105,-7,-104,-172,-151,2,184,210,29,-159,-169,-116,-120,-8,225,186,-104,-43,339,272,-225,-285,114,187,-14,158,477,337,16,45,179,45,-156,-171,-75,31,77,-34,-202,-229,-164,-112,-2,112,34,-119,-49,160,181,4,-106,-8,186,250,115,-8,-1,-61,-202,-102,179,155,-121,-81,239,290,115,159,267,41,-228,-63,287,284,-20,-204,-157,-101,-174,-232,-56,255,328,94,-53,36,11,-217,-228,49,140,-45,-60,109,12,-313,-394,-226,-153,-178,-138,-96,-73,16,11,-215,-365,-244,-130,-145,-76,-21,-204,-296,-6,207,-5,-209,-135,-115,-189,-86,-34,-244,-209,268,447,71,-90,178,183,-131,-134,82,-16,-223,-157,-133,-348,-375,-130,-45,-77,99,201,-86,-292,-7,338,313,117,-46,-220,-281,-96,99,58,-109,-215,-183,-6,125,-24,-241,-108,242,305,42,-131,-13,202,265,149,52,97,127,35,-9,56,57,36,179,300,140,-77,-95,-73,-87,46,211,125,-25,51,150,39,-51,65,170,68,-127,-204,-96,53,96,145,303,322,100,17,194,195,-36,-18,230,190,-114,-226,-86,105,261,236,-21,-195,-152,-181,-259,-17,368,361,41,-120,-67,-9,-6,-78,-192,-174,-20,54,55,143,232,174,56,-12,-31,-25,-94,-263,-259,57,301,220,109,115,43,-34,58,80,-61,3,278,314,123,46,8,-77,3,84,-165,-312,105,468,163,-240,-149,16,-107,-151,49,138,24,-13,76,92,-11,-104,-147,-217,-276,-153,82,98,-75,-58,66,-105,-355,-225,-21,-172,-298,-93,-26,-247,-185,209,309,60,-46,9,-52,-124,-38,49,49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	);
	-- TAMANHO 1060 - Símbolo OFDM parte imaginária, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,-241,-142,-79,-110,-46,-71,-296,-384,-232,-109,17,300,443,217,-3,66,131,-16,-132,-64,31,78,150,181,59,-55,59,201,8,-327,-267,80,90,-225,-240,70,115,-147,-184,64,136,-73,-201,-68,116,121,0,-46,19,12,-155,-341,-401,-342,-250,-197,-172,-110,-78,-175,-203,51,280,108,-189,-172,11,80,137,199,80,-51,88,265,191,87,129,79,-124,-203,-104,-26,-33,-85,-129,-47,129,164,58,44,92,53,53,139,59,-177,-251,-176,-158,-81,88,14,-268,-254,66,195,108,138,211,138,91,111,-100,-466,-465,-32,262,78,-250,-268,-3,153,26,-161,-198,-138,-45,63,35,-146,-126,222,407,129,-168,-117,-36,-211,-380,-298,-89,106,239,191,-11,-91,29,102,24,-58,-112,-179,-112,128,206,-49,-245,-59,190,133,-14,73,212,114,-108,-231,-248,-160,38,128,-31,-134,26,87,-180,-350,-147,-1,-217,-432,-339,-134,-5,125,246,217,47,-112,-151,-115,-150,-249,-210,-77,-146,-270,1,405,262,-189,-178,118,30,-220,-79,180,106,-79,-106,-112,-141,-93,-51,-13,198,425,308,-20,-125,29,162,122,-38,-135,-34,128,186,215,202,4,-107,199,465,137,-321,-258,49,127,67,-36,-198,-147,139,143,-155,-187,-4,-83,-227,-121,-98,-266,-193,34,-35,-163,6,139,66,144,279,76,-185,-129,-73,-194,-162,-40,-181,-347,-180,102,270,382,335,142,165,312,96,-219,-43,238,11,-296,-145,99,97,97,106,-101,-281,-154,1,-66,-142,-47,142,258,89,-318,-436,-27,333,196,-58,-33,86,98,61,-7,-83,-31,102,105,-3,-60,-55,-31,-10,-72,-175,-106,94,120,-28,-69,-15,-49,-51,124,265,197,122,168,114,-152,-357,-266,-73,-69,-142,35,376,419,67,-220,-125,122,213,154,76,51,108,171,117,12,36,128,87,-17,32,175,182,32,-132,-231,-230,-128,-16,67,138,56,-250,-368,3,302,-23,-363,13,511,294,-139,22,371,226,-92,-65,70,9,-45,59,143,127,98,97,136,167,34,-227,-286,-46,137,26,-140,-81,110,140,-56,-232,-165,50,170,133,23,-87,-110,-14,66,45,69,205,223,-28,-320,-322,2,349,374,100,-83,5,79,-58,-176,-73,124,234,216,98,-15,-33,-59,-171,-187,-22,53,-71,-95,90,156,-9,-79,48,69,-82,-88,92,94,-162,-316,-222,-113,-105,-108,-92,-7,200,271,-5,-199,70,278,-47,-332,-62,265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- A saída da convolução vai ter tamanho 1572
	
	component fir_filter 
	generic( 
		Win 		: INTEGER	; -- Input bit width
		Wmult 		: INTEGER	;-- Multiplier bit width 2*W1
		Wadd 		: INTEGER	;-- Adder width = Wmult+log2(L)-1
		Wout 		: INTEGER	;-- Output bit width
		BUTTON_HIGH : STD_LOGIC ;
		LFilter  	: INTEGER	);--Filter Length
	port (
		clk      : in  std_logic	;
		reset    : in  std_logic	;
		i_coeff  : in  ARRAY_COEFF(0 to Lfilter-1)		;
		i_data   : in  std_logic_vector( Win-1 	downto 0)	;
		o_data   : out std_logic_vector( Wout-1 downto 0)   ;
		read_out   : out integer  );
	end component;

	signal i_coeff 	: ARRAY_COEFF(0 to Lfilter-1); 
	signal i_data   : std_logic_vector( Win-1  downto 0);
	signal NOISY	: ARRAY_COEFF(0 to noisy_size-1);

begin
	
	u_fir_filter : fir_filter
	generic map( 
		Win 		 => Win				, -- Input bit width
		Wmult		 => Wmult			,
		Wadd		 => Wadd			,
		Wout 		 => Wout			,-- Output bit width
		BUTTON_HIGH  => BUTTON_HIGH		,
		LFilter  	 => LFilter			) -- Filter length	
	port map(
		clk         => clk       	,
		reset       => reset      	,
		i_coeff     => i_coeff		,
		i_data      => i_data 		,
		o_data     	=> o_data_buffer ,
		read_out  	=> read_out      );

	p_input : process (reset,clk)
		variable control  	: unsigned(11 downto 0):= (others=>'0');
		variable count 		: integer := 0;
		variable count2     : integer := 0;
		variable s			: integer RANGE 0 TO 2**8-1 :=255;
		variable first_time : std_logic := '0';
	begin
		if(reset=BUTTON_HIGH) then
			i_data       <= (others=>'0'); 
			count 		:= 0;
			count2 		:= 0;
			first_time	:='0';
		elsif(rising_edge(clk)) then
			if(first_time='0') then
				for k in 0 to Lfilter-1 loop
					i_coeff(k)  <=  std_logic_vector(to_signed(COEFF_ARRAY(k),Win));
				end loop;			
				for j in 0 to noisy_size-1 loop
					NOISY(j)  <=  std_logic_vector(to_signed(NOISY_ARRAY(j),Win));
				end loop;
				first_time := '1';
			else
				--if(count>=5000 and count<10000) then
				--	s:= 0;
				--elsif (count>=10000) then 
				--	count:=0;
				--	s:=255;
				--end if;
				--i_data<=std_logic_vector(to_unsigned(s,Win));

				--count := count+1;
				--
				--if(count < 5000) then
				--	i_data   <= ('0',others=>'1');
				--elsif(count >= 5000 and count <10000) then
				--	i_data   <= (others=>'0');
				--elsif(count >=10000) then
				--	i_data   <= (others=>'0');
				--	count := 0;
				--end if;				
				--
				-- DELTA, STEP ...........
				--if(control=100 and count2 = 0) then  -- delta
				--	i_data       <= ('0',others=>'1');
				--elsif(control(11)='1' and count2 <3000 ) then  -- step
				--	i_data       <= ('0',others=>'1');
				--	count2 := count2 + 1;
				--else
				--	i_data       <= (others=>'0');
				--end if;
				--control := control + 1;
				------------------------------------------------

				-- DELTA, STEP, STEP, STEP, .......
				--if(control=10) then  -- delta
				--	i_data       <= ('0',others=>'1');
				--elsif(control(7)='1') then  -- step
				--	i_data       <= ('0',others=>'1');
				--else
				--	i_data       <= (others=>'0');
				--end if;
				--control := control + 1;
				-------------------------------------------------
				
				-- NOISY ANALOG SIGNAL
				if(count < noisy_size) then
					i_data <= NOISY(count);
					count := count + 1;
				else
					i_data <= (others=>'0');
				end if;
				-------------------------------------------------

				-- COEFFICIENTS
				if(count < Lfilter-1) then
					o_fir_coeff <= i_coeff(count);
				else
					o_fir_coeff <= (others=>'0');
				end if;
				---------------------------------------------------

				--count := count+1;
			end if;
		end if;
	end process p_input;





end rtl;
